// This holds the blackbox module definitions for the ac97, des3_area, and mc_top

module des3_perf(
output	[63:0]	desOut,
input	[63:0]	desIn,
input	[55:0]	key1,
input	[55:0]	key2,
input	[55:0]	key3,
input		decrypt,
input		clk);
endmodule // des3_perf