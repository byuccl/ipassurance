module potato
   (clk,
    timer_clk,
    reset,
    irq,
    fromhost_data,
    fromhost_updated,
    tohost_data,
    tohost_updated,
    wb_adr_out,
    wb_sel_out,
    wb_cyc_out,
    wb_stb_out,
    wb_we_out,
    wb_dat_out,
    wb_dat_in,
    backdoor,
    wb_ack_in);
  output backdoor;
  input clk;
  input timer_clk;
  input reset;
  input [7:0]irq;
  input [31:0]fromhost_data;
  input fromhost_updated;
  output [31:0]tohost_data;
  output tohost_updated;
  output [31:0]wb_adr_out;
  output [3:0]wb_sel_out;
  output wb_cyc_out;
  output wb_stb_out;
  output wb_we_out;
  output [31:0]wb_dat_out;
  input [31:0]wb_dat_in;
  input wb_ack_in;

  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const0>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const1>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire FSM_sequential_state;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:8]SHIFT_LEFT;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [23:0]SHIFT_RIGHT;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire alu_op;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \alu_op[0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \alu_op[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \alu_op[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \alu_op[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \alu_op[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \alu_op[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire alu_op_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire alu_y_src;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\arbiter/state ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire branch;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \branch[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \branch[2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_28_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_29_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_30_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_31_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_32_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_33_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_34_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_35_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_36_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_37_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_38_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_39_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_40_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_41_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_42_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_43_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_44_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_45_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_46_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_47_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_48_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_49_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_50_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_51_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_52_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_53_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_54_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_55_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_56_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_57_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_58_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_i_59_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_reg_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_reg_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_reg_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_reg_i_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_reg_i_14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_reg_i_15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_reg_i_16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_reg_i_17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_reg_i_18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_reg_i_19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_reg_i_20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_reg_i_21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_reg_i_22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_reg_i_23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_reg_i_24_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_reg_i_25_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_reg_i_26_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_reg_i_27_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_reg_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_reg_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_reg_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_reg_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_reg_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cache_hit_reg_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cancel_fetch_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cl_current_word;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cl_current_word[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cl_current_word[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cl_current_word[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cl_current_word[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cl_load_address;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire clk;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire count_instr_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire count_instr_out_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire count_instruction_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire counter_mtime;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]counter_mtime_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[0]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[0]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[0]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[0]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[12]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[12]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[12]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[12]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[12]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[12]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[12]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[16]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[16]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[16]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[16]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[16]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[16]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[16]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[20]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[20]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[20]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[20]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[20]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[20]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[20]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[24]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[24]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[24]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[24]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[24]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[24]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[24]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[28]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[28]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[28]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[28]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[4]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[4]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[4]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[4]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[4]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[4]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[4]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[8]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[8]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[8]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[8]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[8]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[8]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \counter_mtime_reg[8]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire csr_addr;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_addr[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_addr[10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_addr[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_addr[11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_addr[11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_addr[11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_addr[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_addr[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_addr[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_addr[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_addr[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_addr[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_addr[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_addr[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_addr[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_addr[9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_addr[9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire csr_addr_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire csr_data_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[10]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[10]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[10]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[11]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[11]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[11]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[11]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[13]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[13]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[14]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[14]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[15]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[16]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[16]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[17]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[17]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[18]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[18]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[18]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[19]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[19]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[1]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[1]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[20]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[20]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[21]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[21]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[22]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[22]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[22]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[23]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[23]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[24]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[24]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[25]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[25]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[26]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[26]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[26]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[27]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[27]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[28]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[28]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[29]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[29]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[2]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[2]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[2]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[30]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[30]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[30]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[30]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[30]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[30]_i_5_n_0_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[30]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[30]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[30]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[30]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[31]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[3]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[3]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[3]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[4]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[4]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[4]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[4]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[4]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[4]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[5]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[5]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[6]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[7]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[7]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[8]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out[9]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out_reg[31]_i_17_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out_reg[31]_i_17_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out_reg[31]_i_17_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out_reg[31]_i_22_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out_reg[31]_i_22_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_data_out_reg[31]_i_22_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]csr_read_address_p;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_read_address_p[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_read_address_p[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_read_address_p[0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_read_address_p[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \csr_read_address_p[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire csr_write;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire current_count;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count[0]_i_5__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]current_count_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[0]_i_1__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[0]_i_1__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[0]_i_1__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[0]_i_1__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[0]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[0]_i_1__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[0]_i_1__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[0]_i_1__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[0]_i_1__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[0]_i_1__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[0]_i_1__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[0]_i_1__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[0]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[0]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[0]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[0]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[0]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[0]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[0]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[12]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[12]_i_1__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[12]_i_1__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[12]_i_1__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[12]_i_1__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[12]_i_1__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[12]_i_1__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[12]_i_1__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[12]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[12]_i_1__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[12]_i_1__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[12]_i_1__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[12]_i_1__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[12]_i_1__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[12]_i_1__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[12]_i_1__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[12]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[12]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[12]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[12]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[12]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[12]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[12]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[16]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[16]_i_1__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[16]_i_1__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[16]_i_1__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[16]_i_1__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[16]_i_1__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[16]_i_1__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[16]_i_1__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[16]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[16]_i_1__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[16]_i_1__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[16]_i_1__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[16]_i_1__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[16]_i_1__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[16]_i_1__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[16]_i_1__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[16]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[16]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[16]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[16]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[16]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[16]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[16]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[20]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[20]_i_1__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[20]_i_1__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[20]_i_1__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[20]_i_1__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[20]_i_1__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[20]_i_1__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[20]_i_1__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[20]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[20]_i_1__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[20]_i_1__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[20]_i_1__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[20]_i_1__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[20]_i_1__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[20]_i_1__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[20]_i_1__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[20]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[20]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[20]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[20]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[20]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[20]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[20]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[24]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[24]_i_1__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[24]_i_1__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[24]_i_1__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[24]_i_1__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[24]_i_1__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[24]_i_1__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[24]_i_1__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[24]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[24]_i_1__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[24]_i_1__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[24]_i_1__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[24]_i_1__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[24]_i_1__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[24]_i_1__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[24]_i_1__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[24]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[24]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[24]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[24]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[24]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[24]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[24]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[28]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[28]_i_1__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[28]_i_1__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[28]_i_1__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[28]_i_1__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[28]_i_1__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[28]_i_1__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[28]_i_1__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[28]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[28]_i_1__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[28]_i_1__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[28]_i_1__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[28]_i_1__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[28]_i_1__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[28]_i_1__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[28]_i_1__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[28]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[28]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[28]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[28]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[28]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[28]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[28]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[32]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[32]_i_1__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[32]_i_1__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[32]_i_1__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[32]_i_1__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[32]_i_1__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[32]_i_1__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[32]_i_1__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[32]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[32]_i_1__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[32]_i_1__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[32]_i_1__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[32]_i_1__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[32]_i_1__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[32]_i_1__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[32]_i_1__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[32]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[32]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[32]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[32]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[32]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[32]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[32]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[32]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[36]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[36]_i_1__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[36]_i_1__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[36]_i_1__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[36]_i_1__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[36]_i_1__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[36]_i_1__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[36]_i_1__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[36]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[36]_i_1__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[36]_i_1__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[36]_i_1__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[36]_i_1__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[36]_i_1__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[36]_i_1__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[36]_i_1__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[36]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[36]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[36]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[36]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[36]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[36]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[36]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[36]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[40]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[40]_i_1__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[40]_i_1__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[40]_i_1__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[40]_i_1__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[40]_i_1__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[40]_i_1__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[40]_i_1__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[40]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[40]_i_1__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[40]_i_1__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[40]_i_1__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[40]_i_1__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[40]_i_1__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[40]_i_1__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[40]_i_1__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[40]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[40]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[40]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[40]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[40]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[40]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[40]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[40]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[44]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[44]_i_1__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[44]_i_1__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[44]_i_1__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[44]_i_1__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[44]_i_1__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[44]_i_1__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[44]_i_1__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[44]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[44]_i_1__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[44]_i_1__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[44]_i_1__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[44]_i_1__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[44]_i_1__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[44]_i_1__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[44]_i_1__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[44]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[44]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[44]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[44]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[44]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[44]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[44]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[44]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[48]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[48]_i_1__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[48]_i_1__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[48]_i_1__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[48]_i_1__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[48]_i_1__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[48]_i_1__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[48]_i_1__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[48]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[48]_i_1__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[48]_i_1__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[48]_i_1__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[48]_i_1__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[48]_i_1__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[48]_i_1__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[48]_i_1__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[48]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[48]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[48]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[48]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[48]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[48]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[48]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[48]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[4]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[4]_i_1__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[4]_i_1__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[4]_i_1__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[4]_i_1__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[4]_i_1__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[4]_i_1__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[4]_i_1__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[4]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[4]_i_1__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[4]_i_1__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[4]_i_1__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[4]_i_1__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[4]_i_1__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[4]_i_1__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[4]_i_1__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[4]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[4]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[4]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[4]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[4]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[4]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[4]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[52]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[52]_i_1__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[52]_i_1__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[52]_i_1__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[52]_i_1__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[52]_i_1__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[52]_i_1__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[52]_i_1__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[52]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[52]_i_1__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[52]_i_1__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[52]_i_1__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[52]_i_1__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[52]_i_1__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[52]_i_1__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[52]_i_1__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[52]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[52]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[52]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[52]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[52]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[52]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[52]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[52]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[56]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[56]_i_1__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[56]_i_1__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[56]_i_1__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[56]_i_1__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[56]_i_1__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[56]_i_1__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[56]_i_1__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[56]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[56]_i_1__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[56]_i_1__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[56]_i_1__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[56]_i_1__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[56]_i_1__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[56]_i_1__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[56]_i_1__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[56]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[56]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[56]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[56]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[56]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[56]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[56]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[56]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[60]_i_1__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[60]_i_1__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[60]_i_1__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[60]_i_1__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[60]_i_1__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[60]_i_1__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[60]_i_1__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[60]_i_1__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[60]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[60]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[60]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[60]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[8]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[8]_i_1__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[8]_i_1__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[8]_i_1__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[8]_i_1__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[8]_i_1__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[8]_i_1__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[8]_i_1__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[8]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[8]_i_1__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[8]_i_1__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[8]_i_1__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[8]_i_1__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[8]_i_1__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[8]_i_1__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[8]_i_1__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[8]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[8]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[8]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[8]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[8]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[8]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \current_count_reg[8]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:25]data0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]data12;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]data14;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]data16;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]data8;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire decode_exception_cause;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire decode_exception_cause1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \decode_exception_cause[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \decode_exception_cause[0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \decode_exception_cause[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \decode_exception_cause[0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \decode_exception_cause[0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \decode_exception_cause[0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \decode_exception_cause[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \decode_exception_cause[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \decode_exception_cause[2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \decode_exception_cause[2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \decode_exception_cause[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \decode_exception_cause[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \decode_exception_cause[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire decode_exception_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire decode_exception_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire decode_exception_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire decode_exception_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire decode_exception_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire decode_exception_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]dmem_address;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:2]dmem_address__0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]dmem_address_p;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_address_p[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_address_p[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:8]dmem_data_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire dmem_data_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[23]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[23]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[23]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[26]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[30]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out[9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]dmem_data_out_p;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out_p[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out_p[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out_p[31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out_p[31]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out_p[31]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_data_out_p[31]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/dmem_data_out_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/state ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/state[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/state_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if/state_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire dmem_if_inputs;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire dmem_if_outputs;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\dmem_if_outputs[adr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\dmem_if_outputs[dat] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\dmem_if_outputs[sel] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dmem_if_outputs[we] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire dmem_r_ack_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire dmem_read_ack;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire dmem_write_ack;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire dmem_write_req;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire exception_context_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][16]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][17]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][18]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][19]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][1]_i_3_n_0_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][20]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][21]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][22]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][23]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][24]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][25]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][26]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][27]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][28]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][29]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][30]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][31]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][31]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[badaddr][9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][0]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][0]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][0]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][0]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][0]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][0]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][0]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][0]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][2]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][2]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][5]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][5]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][5]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][5]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][5]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[cause][5]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[ie1]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[ie1]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[ie1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[ie1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[ie1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[ie1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[ie1]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[ie1]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[ie1]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[ie]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \exception_context_out[ie]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]fromhost;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]fromhost_data;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire fromhost_updated;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/cache_hit ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/cache_hit0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/cache_memory_reg_0_n_51 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/cache_memory_reg_0_n_52 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/cache_memory_reg_0_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/cache_memory_reg_0_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/cache_memory_reg_0_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/cache_memory_reg_0_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/cache_memory_reg_1_n_27 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/cache_memory_reg_1_n_28 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/cache_memory_reg_1_n_53 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/cache_memory_reg_1_n_54 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/cache_memory_reg_1_n_55 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/cache_memory_reg_1_n_56 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/cache_memory_reg_1_n_57 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/cache_memory_reg_1_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/cache_memory_reg_1_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/cache_memory_reg_1_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/cl_current_word_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/cl_current_word_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/cl_current_word_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:4]\icache/cl_load_address ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [125:0]\icache/current_cache_line ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\icache/input_address_word ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/input_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/input_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/input_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/input_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/input_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/input_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/input_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]\icache/load_buffer ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/p_1_in10_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/p_3_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/read_ack ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/state_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/state_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/state_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/store_cache_line__1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/store_cache_line_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_0_63_0_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_0_63_0_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_0_63_0_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_0_63_12_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_0_63_12_14_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_0_63_12_14_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_0_63_15_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_0_63_15_17_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_0_63_15_17_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_0_63_18_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_0_63_18_20_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_0_63_18_20_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_0_63_3_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_0_63_3_5_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_0_63_3_5_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_0_63_6_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_0_63_6_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_0_63_6_8_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_0_63_9_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_0_63_9_11_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_0_63_9_11_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_64_127_0_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_64_127_0_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_64_127_0_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_64_127_12_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_64_127_12_14_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_64_127_12_14_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_64_127_15_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_64_127_15_17_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_64_127_15_17_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_64_127_18_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_64_127_18_20_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_64_127_18_20_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_64_127_3_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_64_127_3_5_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_64_127_3_5_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_64_127_6_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_64_127_6_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_64_127_6_8_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_64_127_9_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_64_127_9_11_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/tag_memory_reg_64_127_9_11_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache/to_std_logic ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]\icache/valid ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire icache_inputs;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire icache_outputs;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:2]\icache_outputs[adr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache_outputs[sel] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \icache_outputs[stb] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ie1_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ie1_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ie_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ie_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ie_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ie_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ie_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire imem_ack;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:2]imem_address;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:2]imem_data;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire immediate;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[13]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[14]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[16]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[16]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[17]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[17]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[18]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[18]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[19]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[19]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[30]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[30]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[30]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \immediate[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire input_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire input_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire input_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire input_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire input_carry__0_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire input_carry__0_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire input_carry__0_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire input_carry__0_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire input_carry__0_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire input_carry_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire input_carry_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire input_carry_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire input_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire input_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire input_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire input_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire input_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire input_carry_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire input_carry_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire input_carry_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire input_carry_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire instruction;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]irq;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire load_buffer;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[101]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[102]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[103]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[104]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[105]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[106]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[107]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[108]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[109]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[110]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[111]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[112]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[113]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[114]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[115]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[116]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[117]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[118]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[119]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[120]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[121]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[122]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[123]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[124]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[125]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[126]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[127]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[127]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[127]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[63]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[64]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[65]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[66]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[67]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[68]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[69]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[70]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[71]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[72]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[73]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[74]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[75]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[76]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[77]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[78]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[79]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[80]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[81]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[82]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[83]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[84]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[85]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[86]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[87]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[88]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[89]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[90]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[91]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[92]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[93]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[94]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[95]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[95]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[96]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[97]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[98]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \load_buffer[99]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]mbadaddr;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mbadaddr[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire mem_op;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_100_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_101_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_102_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_103_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_104_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_105_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_106_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_107_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_108_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_109_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_110_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_111_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_112_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_114_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_115_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_116_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_117_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_118_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_119_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_120_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_121_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_123_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_124_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_125_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_126_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_127_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_128_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_129_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_130_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_132_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_133_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_134_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_135_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_136_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_137_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_138_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_139_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_141_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_142_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_143_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_144_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_145_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_146_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_147_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_148_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_149_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_150_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_151_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_152_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_153_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_154_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_155_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_156_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_157_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_158_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_159_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_160_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_161_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_162_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_163_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_164_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_165_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_166_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_167_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_168_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_169_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_170_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_171_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_172_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_173_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_174_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_175_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_176_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_177_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_178_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_179_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_180_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_52_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_53_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_54_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_55_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_57_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_58_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_60_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_61_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_62_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_63_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_65_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_66_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_67_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_68_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_70_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_71_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_72_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_73_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_74_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_75_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_76_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_77_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_79_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_80_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_81_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_82_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_83_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_84_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_85_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_86_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_88_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_89_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_90_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_91_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_92_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_93_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_94_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_95_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_97_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_98_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op[2]_i_99_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]mem_op_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_11_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_11_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_11_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_122_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_122_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_122_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_122_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_12_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_12_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_12_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_131_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_131_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_131_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_131_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_13_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_13_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_13_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_140_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_140_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_140_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_140_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_14_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_14_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_14_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_15_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_15_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_15_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_19_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_19_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_19_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_23_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_23_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_23_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_32_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_32_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_41_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_41_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_41_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_50_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_50_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_50_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_59_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_59_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_59_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_59_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_64_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_64_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_64_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_64_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_69_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_69_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_69_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_69_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_78_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_78_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_78_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_78_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_87_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_87_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_87_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_87_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_96_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_96_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_96_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_96_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_9_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_op_reg[2]_i_9_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]mem_size;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_size[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_size[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_size[0]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_size[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_size[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_size[1]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_size[1]_repN_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mem_size[1]_repN_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]mepc;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mepc[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mepc[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire mie;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mie[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]mscratch;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mscratch[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]mtime_compare;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtime_compare[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtime_compare[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtime_compare[31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]mtvec;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire mtvec_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[18]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[22]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[26]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[30]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mtvec_out[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_0_in0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_0_in0_repN;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]p_0_out1_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_1_in0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]p_1_out0_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]p_1_out2_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]p_2_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]pc;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[11]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[11]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[11]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[15]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[15]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[15]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[16]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[17]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[18]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[19]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[19]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[19]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[19]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[19]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[20]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[21]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[22]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[23]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[23]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[23]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[23]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[23]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[24]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[25]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[26]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[27]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[27]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[27]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[27]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[27]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[28]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[29]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[30]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[31]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[31]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[31]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[31]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[31]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[4]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[7]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[7]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[7]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]pc_next;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]pc_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[11]_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[11]_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[11]_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[11]_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[12]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[12]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[12]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[12]_i_4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[12]_i_4_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[12]_i_4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[12]_i_4_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[12]_i_4_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[12]_i_4_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[12]_i_4_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[15]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[15]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[15]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[15]_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[15]_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[15]_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[15]_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[16]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[16]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[16]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[16]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[16]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[16]_i_4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[16]_i_4_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[16]_i_4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[16]_i_4_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[16]_i_4_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[16]_i_4_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[16]_i_4_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[19]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[19]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[19]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[19]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[19]_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[19]_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[19]_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[19]_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[20]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[20]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[20]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[20]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[20]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[20]_i_4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[20]_i_4_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[20]_i_4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[20]_i_4_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[20]_i_4_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[20]_i_4_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[20]_i_4_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[23]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[23]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[23]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[23]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[23]_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[23]_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[23]_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[23]_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[24]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[24]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[24]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[24]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[24]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[24]_i_4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[24]_i_4_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[24]_i_4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[24]_i_4_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[24]_i_4_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[24]_i_4_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[24]_i_4_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[27]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[27]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[27]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[27]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[27]_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[27]_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[27]_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[27]_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[28]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[28]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[28]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[28]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[28]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[28]_i_4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[28]_i_4_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[28]_i_4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[28]_i_4_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[28]_i_4_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[28]_i_4_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[28]_i_4_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[31]_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[31]_i_5_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[31]_i_5_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[31]_i_5_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[31]_i_5_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[31]_i_9_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[31]_i_9_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[31]_i_9_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[31]_i_9_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[3]_i_4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[3]_i_4_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[3]_i_4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[3]_i_4_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[3]_i_4_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[3]_i_4_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[3]_i_4_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[4]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[4]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[4]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[4]_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[4]_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[4]_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[4]_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[7]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[7]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[7]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[7]_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[7]_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[7]_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[7]_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[8]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[8]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[8]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[8]_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[8]_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[8]_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[8]_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/csr_read_data ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_read_writeable ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/csr_unit/counter_mtime_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/cycle_counter/current_count_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/ie1__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/ie__7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/instret_counter/current_count_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/mscratch__4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/mtime_compare__4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/mtvec_out1__6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/read_data_out2__3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/read_data_out2_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/read_data_out2_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/read_data_out2_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/csr_unit/read_data_out__582 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/software_interrupt__5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_counter/current_count_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_interrupt0__8 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_interrupt0_inferred__0_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_interrupt0_inferred__0_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_interrupt0_inferred__0_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_interrupt0_inferred__0_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_interrupt0_inferred__0_carry__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_interrupt0_inferred__0_carry__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_interrupt0_inferred__0_carry__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_interrupt0_inferred__0_carry__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_interrupt0_inferred__0_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_interrupt0_inferred__0_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_interrupt0_inferred__0_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/timer_interrupt0_inferred__0_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/tohost_data0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/csr_unit/tohost_data1__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [9:0]\processor/decode/csr_addr__40 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/decode/instruction_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/decode/instruction_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/decode/instruction_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/decode/instruction_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/decode/instruction_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\processor/dmem_data_size_p ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/dmem_read_req_p ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/dmem_write_req_p ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\processor/ex_branch ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/ex_count_instruction ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\processor/ex_csr_address ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/ex_csr_address[3]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/ex_csr_address[6]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/ex_csr_address[6]_repN_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/ex_csr_address[7]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\processor/ex_csr_write ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/ex_dmem_data_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\processor/ex_dmem_data_size ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/ex_dmem_read_req ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/ex_dmem_write_req ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/ex_exception_context ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/ex_exception_context[badaddr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:0]\processor/ex_exception_context[cause] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/ex_exception_context[ie] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\processor/ex_mem_op ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/ex_mem_size ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/ex_pc ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\processor/ex_rd_address ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/ex_rd_data ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/ex_rd_write ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/exception_target ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/execute/alu_instance/data3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/execute/alu_instance/data4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/execute/alu_instance/data5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/execute/alu_instance/data6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\processor/execute/alu_instance/data7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:1]\processor/execute/alu_instance/data9 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\processor/execute/alu_op ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/execute/alu_x ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/execute/alu_x[27]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:1]\processor/execute/alu_x_mux/data3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\processor/execute/alu_x_src ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/execute/alu_y ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:1]\processor/execute/alu_y_mux/data3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\processor/execute/alu_y_src ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/execute/branch_comparator/data0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/execute/branch_comparator/data1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/execute/branch_comparator/data2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/execute/branch_comparator/data3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/execute/branch_comparator/data4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/execute/branch_comparator/data5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/execute/branch_condition ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/execute/csr_alu_instance/b ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/execute/csr_value_forwarded3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/execute/csr_value_forwarded30_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/execute/csr_writeable ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/execute/decode_exception ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\processor/execute/decode_exception_cause ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/execute/exception_taken0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\processor/execute/funct3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/execute/immediate ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:3]\processor/execute/mie ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/execute/mtvec ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:5]\processor/execute/mtvec_forwarded ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/execute/rd_write_out0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\processor/execute/rs1_addr ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/execute/rs1_addr[0]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/execute/rs1_forwarded ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/execute/rs1_forwarded[7]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\processor/execute/rs2_addr ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\processor/execute/shamt ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/fetch/cancel_fetch ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\processor/id_alu_op ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\processor/id_alu_x_src ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\processor/id_alu_y_src ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\processor/id_branch ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/id_count_instruction ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/id_csr_use_immediate ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\processor/id_csr_write ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/id_exception ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\processor/id_exception_cause ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\processor/id_funct3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/id_immediate ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\processor/id_mem_op ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/id_mem_size ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/id_pc ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\processor/id_rd_address ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/id_rd_write ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\processor/id_rs1_address ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\processor/id_shamt ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/ie ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/ie1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\processor/mem_csr_address ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/mem_csr_address[4]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/mem_csr_address[4]_repN_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/mem_csr_data ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\processor/mem_csr_write ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/mem_exception ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/mem_exception_context ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/mem_exception_context[badaddr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:0]\processor/mem_exception_context[cause] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/mem_exception_context[ie] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\processor/mem_mem_op ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/mem_mem_op[1]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/mem_mem_op[1]_repN_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/mem_mem_op[1]_repN_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\processor/mem_rd_address ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/mem_rd_data ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/mem_rd_data[7]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/mem_rd_data[7]_repN_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/mem_rd_write ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/memory/csr_write_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/memory/csr_write_out[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/memory/exception_out0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/memory/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/mie ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/mtvec ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/regfile/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\processor/rs1_address ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\processor/rs1_address_p ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/rs1_data ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\processor/rs2_address ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\processor/rs2_address_p ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/rs2_data ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/software_interrupt ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/timer_interrupt ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\processor/wb_csr_address ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/wb_csr_data ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\processor/wb_csr_write ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/wb_exception ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/wb_exception_context ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/wb_exception_context[badaddr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:0]\processor/wb_exception_context[cause] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/wb_exception_context[ie] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\processor/wb_rd_address ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\processor/wb_rd_data ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/wb_rd_write ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \processor/writeback/count_instr_out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]rd_data;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_52_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_54_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_55_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_57_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_58_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_59_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_60_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_61_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_62_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_63_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_64_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_65_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_66_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_67_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_68_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_69_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[10]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[10]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[10]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[10]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[10]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[10]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[10]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[10]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[10]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[10]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[10]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[11]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[12]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[12]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[12]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[12]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[12]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[12]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[12]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[13]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[13]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[13]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[13]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[13]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[13]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[13]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[13]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[13]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[13]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[14]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[14]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[14]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[14]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[14]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[14]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[14]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[14]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[14]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[14]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[15]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[16]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[16]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[16]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[16]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[16]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[16]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[16]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[16]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[16]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[16]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[16]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[16]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[17]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[17]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[17]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[17]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[17]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[17]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[17]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[17]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[17]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[17]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[17]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[17]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[18]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[18]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[18]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[18]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[18]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[18]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[18]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[18]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[18]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[18]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[18]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[18]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[19]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[1]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[1]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[1]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[1]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[1]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[20]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[20]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[20]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[20]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[20]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[20]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[20]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[20]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[20]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[20]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[20]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[20]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[21]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[21]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[21]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[21]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[21]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[21]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[21]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[21]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[21]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[21]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[21]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[21]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[22]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[22]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[22]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[22]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[22]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[22]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[22]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[22]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[22]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[22]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[22]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[22]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[23]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[24]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[24]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[24]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[24]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[24]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[24]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[24]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[24]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[24]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[24]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[24]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[25]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[25]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[25]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[25]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[25]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[25]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[25]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[25]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[25]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[25]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[25]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[26]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[26]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[26]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[26]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[26]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[26]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[26]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[26]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[26]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[26]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[26]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[27]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[28]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[28]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[28]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[28]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[28]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[28]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[28]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[28]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[28]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[28]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[28]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[29]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[29]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[29]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[29]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[29]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[29]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[29]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[29]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[29]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[2]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[2]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[2]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[2]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[2]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[2]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[2]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[30]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[31]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[31]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[31]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[31]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[31]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[31]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[31]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[31]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[31]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[31]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[31]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[31]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[31]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[31]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[31]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[31]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[31]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[31]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[31]_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[31]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[31]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[3]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[3]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[3]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[3]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[3]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[3]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[3]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[3]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[3]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[3]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[3]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[3]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[3]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[3]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[3]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[3]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[3]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[4]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[4]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[4]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[4]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[4]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[4]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[4]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[4]_i_8_n_0_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[5]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[5]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[5]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[5]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[5]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[5]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[5]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[6]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[6]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[6]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[6]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[6]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[6]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[6]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[7]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[8]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[8]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[8]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[8]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[8]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[8]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[8]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[9]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[9]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[9]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[9]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[9]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[9]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[9]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[9]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data[9]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_data_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_out[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_out[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_out[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_out[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_out[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_out[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_out[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_out[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_out[31]_i_2_n_0_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_out[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_out[31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_out[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_out[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]rd_data_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_22_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_22_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_22_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_30_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_30_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_30_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_39_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_39_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_39_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_44_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_44_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_44_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_53_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_53_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_53_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_53_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_9_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_9_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[0]_i_9_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[11]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[11]_i_12_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[11]_i_12_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[11]_i_12_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[11]_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[11]_i_40_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[11]_i_40_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[11]_i_40_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[11]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[11]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[11]_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[11]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[12]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[12]_i_14_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[12]_i_14_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[12]_i_14_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[15]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[15]_i_12_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[15]_i_12_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[15]_i_12_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[15]_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[15]_i_39_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[15]_i_39_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[15]_i_39_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[15]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[15]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[15]_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[15]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[16]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[16]_i_15_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[16]_i_15_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[16]_i_15_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[19]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[19]_i_13_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[19]_i_13_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[19]_i_13_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[19]_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[19]_i_41_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[19]_i_41_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[19]_i_41_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[19]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[19]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[19]_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[19]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[20]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[20]_i_15_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[20]_i_15_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[20]_i_15_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[23]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[23]_i_12_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[23]_i_12_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[23]_i_12_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[23]_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[23]_i_39_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[23]_i_39_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[23]_i_39_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[23]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[23]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[23]_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[23]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[24]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[24]_i_14_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[24]_i_14_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[24]_i_14_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[27]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[27]_i_13_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[27]_i_13_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[27]_i_13_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[27]_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[27]_i_40_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[27]_i_40_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[27]_i_40_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[27]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[27]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[27]_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[27]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[2]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[2]_i_11_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[2]_i_11_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[2]_i_11_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[2]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[2]_i_13_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[2]_i_13_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[2]_i_13_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[31]_i_15_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[31]_i_17_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[31]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[31]_i_32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[31]_i_32_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[31]_i_32_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[31]_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[31]_i_36_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[31]_i_36_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[31]_i_36_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[3]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[3]_i_12_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[3]_i_12_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[3]_i_12_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[3]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[3]_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[3]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[7]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[7]_i_12_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[7]_i_12_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[7]_i_12_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[7]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[7]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[7]_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[7]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[8]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[8]_i_14_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[8]_i_14_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rd_data_reg[8]_i_14_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_write_out_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire read_ack_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire read_data_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire read_data_out2_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire read_data_out2_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire read_data_out2_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire read_data_out2_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[10]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[10]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[10]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[10]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[11]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[11]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[11]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[12]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[12]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[13]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[13]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[13]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[13]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[14]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[14]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[14]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[14]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[15]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[15]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[15]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[16]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[16]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[16]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[16]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[17]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[17]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[17]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[17]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[18]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[18]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[18]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[18]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[18]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[19]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[19]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[19]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[19]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[1]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[20]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[20]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[20]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[20]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[21]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[21]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[21]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[21]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[22]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[22]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[22]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[22]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[22]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[23]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[23]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[23]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[23]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[24]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[24]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[24]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[24]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[25]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[25]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[25]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[25]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[26]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[26]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[26]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[26]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[26]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[27]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[27]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[27]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[27]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[28]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[28]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[28]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[28]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[29]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[29]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[29]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[29]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[2]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[30]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[30]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[30]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[30]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[30]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[31]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[4]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[4]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[5]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[5]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[5]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[6]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[6]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[6]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[7]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[7]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[7]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[8]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[8]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[9]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[9]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out[9]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire read_data_out_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[10]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[13]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[14]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[16]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[17]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[18]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[19]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[20]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[21]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[22]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[23]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[24]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[25]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[26]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[27]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[28]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[29]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[30]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[31]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[5]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[6]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \read_data_out_reg[9]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire registers_reg_r1_0_31_0_5_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire registers_reg_r1_0_31_0_5_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire registers_reg_r1_0_31_0_5_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire registers_reg_r1_0_31_0_5_i_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire registers_reg_r1_0_31_0_5_i_14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire registers_reg_r1_0_31_0_5_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire registers_reg_r1_0_31_0_5_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire reset;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rs1_data;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rs1_data[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rs2_data;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rs2_data[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire software_interrupt_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire state;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \state[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \state[1]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \state[1]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \state[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \state[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire store_cache_line_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire tag_memory_reg_0_63_0_2_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire tag_memory_reg_0_63_0_2_i_15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire tag_memory_reg_0_63_0_2_i_16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire tag_memory_reg_0_63_0_2_i_18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire tag_memory_reg_0_63_0_2_i_19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire tag_memory_reg_0_63_0_2_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire tag_memory_reg_0_63_0_2_i_20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire tag_memory_reg_0_63_0_2_i_21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire tag_memory_reg_0_63_0_2_i_22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire tag_memory_reg_0_63_0_2_i_23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire tag_memory_reg_0_63_0_2_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire tag_memory_reg_0_63_0_2_i_8_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire tag_memory_reg_0_63_0_2_i_8_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire tag_memory_reg_0_63_0_2_i_8_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire tag_memory_reg_0_63_0_2_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire tag_memory_reg_64_127_0_2_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire timer_clk;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire timer_interrupt0_inferred__0_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire timer_interrupt0_inferred__0_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire timer_interrupt0_inferred__0_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire timer_interrupt0_inferred__0_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire timer_interrupt0_inferred__0_carry__1_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire timer_interrupt0_inferred__0_carry__1_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire timer_interrupt0_inferred__0_carry__1_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire timer_interrupt0_inferred__0_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire timer_interrupt0_inferred__0_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire timer_interrupt0_inferred__0_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire timer_interrupt0_inferred__0_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire timer_interrupt_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire timer_interrupt_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire timer_interrupt_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]tohost_data;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tohost_data[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tohost_data[31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tohost_data[31]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire tohost_updated;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire valid;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[100]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[101]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[102]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[103]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[104]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[105]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[106]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[107]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[108]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[109]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[110]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[111]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[111]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[112]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[112]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[113]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[113]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[114]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[114]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[115]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[115]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[116]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[116]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[117]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[117]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[118]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[118]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[119]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[119]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[120]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[120]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[121]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[121]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[122]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[122]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[123]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[123]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[124]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[124]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[125]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[125]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[126]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[126]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[127]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[127]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[127]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[18]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[22]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[26]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[30]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[32]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[33]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[34]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[35]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[36]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[37]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[38]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[39]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[40]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[41]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[42]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[43]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[44]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[45]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[46]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[47]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[47]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[48]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[49]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[50]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[51]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[52]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[53]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[54]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[55]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[56]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[57]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[58]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[59]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[60]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[61]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[62]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[63]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[63]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[64]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[65]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[66]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[67]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[68]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[69]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[70]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[71]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[72]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[73]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[74]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[75]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[76]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[77]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[78]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[79]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[79]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[80]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[81]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[82]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[83]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[84]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[85]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[86]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[87]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[88]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[89]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[90]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[91]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[92]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[93]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[94]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[95]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[95]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[96]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[97]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[98]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[99]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \valid[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire wb_ack_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]wb_adr_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire wb_cyc_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]wb_dat_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]wb_dat_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire wb_outputs;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][12]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][13]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][15]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][16]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][18]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][19]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][21]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][22]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][24]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][25]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][26]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][27]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][28]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][2]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][30]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][31]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][31]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][3]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][6]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][7]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[adr][9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[cyc]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[cyc]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[cyc]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[cyc]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][24]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][24]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][25]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][25]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][26]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][26]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][27]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][27]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][28]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][28]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][29]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][29]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][30]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][30]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[dat][7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[sel][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[sel][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[sel][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[sel][3]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[sel][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[stb]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[we]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \wb_outputs[we]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]wb_sel_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire wb_stb_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire wb_we_out;

  assign backdoor =  wb_we_out ;

  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD850)) 
    \FSM_sequential_state[0]_i_1 
       (.I0(\arbiter/state [1]),
        .I1(\arbiter/state [0]),
        .I2(icache_outputs),
        .I3(dmem_if_outputs),
        .O(FSM_sequential_state));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hAB00)) 
    \FSM_sequential_state[1]_i_1 
       (.I0(\arbiter/state [1]),
        .I1(\arbiter/state [0]),
        .I2(icache_outputs),
        .I3(dmem_if_outputs),
        .O(\FSM_sequential_state[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND
       (.G(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC
       (.P(\<const1>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFEE7)) 
    \alu_op[0]_i_1 
       (.I0(\processor/decode/instruction_reg_n_0_ ),
        .I1(\processor/decode/instruction_reg_n_0_[3] ),
        .I2(\processor/decode/instruction_reg_n_0_[4] ),
        .I3(\processor/decode/instruction_reg_n_0_[6] ),
        .I4(alu_op_reg),
        .O(\processor/id_alu_op [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h11415555)) 
    \alu_op[0]_i_3 
       (.I0(\processor/decode/instruction_reg_n_0_[3] ),
        .I1(\processor/id_funct3 [0]),
        .I2(\processor/id_csr_use_immediate ),
        .I3(\processor/id_funct3 [1]),
        .I4(\processor/decode/instruction_reg_n_0_[4] ),
        .O(alu_op));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBEBBBEBAAAAAAAAA)) 
    \alu_op[0]_i_4 
       (.I0(\processor/decode/instruction_reg_n_0_[3] ),
        .I1(\processor/id_funct3 [0]),
        .I2(\processor/id_funct3 [1]),
        .I3(\processor/id_csr_use_immediate ),
        .I4(\alu_op[3]_i_3_n_0 ),
        .I5(\processor/decode/instruction_reg_n_0_[4] ),
        .O(\alu_op[0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF7FFF7FBB6E8A6E)) 
    \alu_op[1]_i_1 
       (.I0(\processor/decode/instruction_reg_n_0_[6] ),
        .I1(\processor/decode/instruction_reg_n_0_ ),
        .I2(\processor/decode/instruction_reg_n_0_[5] ),
        .I3(\processor/decode/instruction_reg_n_0_[4] ),
        .I4(\alu_op[1]_i_2_n_0 ),
        .I5(\processor/decode/instruction_reg_n_0_[3] ),
        .O(\processor/id_alu_op [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000046074606)) 
    \alu_op[1]_i_2 
       (.I0(\processor/id_funct3 [1]),
        .I1(\processor/id_csr_use_immediate ),
        .I2(\processor/id_funct3 [0]),
        .I3(\alu_op[3]_i_3_n_0 ),
        .I4(\processor/decode/instruction_reg_n_0_[5] ),
        .I5(\processor/decode/instruction_reg_n_0_[6] ),
        .O(\alu_op[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0A0000000AA0F0CF)) 
    \alu_op[2]_i_1 
       (.I0(\processor/decode/instruction_reg_n_0_[5] ),
        .I1(\alu_op[2]_i_2_n_0 ),
        .I2(\processor/decode/instruction_reg_n_0_[4] ),
        .I3(\processor/decode/instruction_reg_n_0_ ),
        .I4(\processor/decode/instruction_reg_n_0_[6] ),
        .I5(\processor/decode/instruction_reg_n_0_[3] ),
        .O(\processor/id_alu_op [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h08C3)) 
    \alu_op[2]_i_2 
       (.I0(\alu_op[3]_i_3_n_0 ),
        .I1(\processor/id_funct3 [0]),
        .I2(\processor/id_funct3 [1]),
        .I3(\processor/id_csr_use_immediate ),
        .O(\alu_op[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF7FFF7FFF6E026E)) 
    \alu_op[3]_i_1 
       (.I0(\processor/decode/instruction_reg_n_0_[6] ),
        .I1(\processor/decode/instruction_reg_n_0_ ),
        .I2(\processor/decode/instruction_reg_n_0_[5] ),
        .I3(\processor/decode/instruction_reg_n_0_[4] ),
        .I4(\alu_op[3]_i_2_n_0 ),
        .I5(\processor/decode/instruction_reg_n_0_[3] ),
        .O(\processor/id_alu_op [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA00000444)) 
    \alu_op[3]_i_2 
       (.I0(\processor/decode/instruction_reg_n_0_ ),
        .I1(\processor/id_funct3 [0]),
        .I2(\alu_op[3]_i_3_n_0 ),
        .I3(\processor/id_csr_use_immediate ),
        .I4(\processor/id_funct3 [1]),
        .I5(\processor/decode/instruction_reg_n_0_[6] ),
        .O(\alu_op[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \alu_op[3]_i_3 
       (.I0(\alu_op[3]_i_4_n_0 ),
        .I1(data0[26]),
        .I2(data0[25]),
        .I3(data0[28]),
        .I4(data0[27]),
        .O(\alu_op[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \alu_op[3]_i_4 
       (.I0(data0[30]),
        .I1(data0[29]),
        .I2(data0[31]),
        .O(\alu_op[3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \alu_op_reg[0]_i_2 
       (.I0(alu_op),
        .I1(\alu_op[0]_i_4_n_0 ),
        .O(alu_op_reg),
        .S(\processor/decode/instruction_reg_n_0_[5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair52" *) 
  LUT5 #(
    .INIT(32'h01200020)) 
    \alu_x_src[0]_i_1 
       (.I0(\processor/decode/instruction_reg_n_0_ ),
        .I1(\processor/decode/instruction_reg_n_0_[3] ),
        .I2(\processor/decode/instruction_reg_n_0_[4] ),
        .I3(\processor/decode/instruction_reg_n_0_[6] ),
        .I4(\processor/decode/instruction_reg_n_0_[5] ),
        .O(\processor/id_alu_x_src [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00044000)) 
    \alu_x_src[1]_i_1 
       (.I0(\processor/decode/instruction_reg_n_0_[3] ),
        .I1(\processor/decode/instruction_reg_n_0_[4] ),
        .I2(\processor/decode/instruction_reg_n_0_[5] ),
        .I3(\processor/decode/instruction_reg_n_0_[6] ),
        .I4(\processor/decode/instruction_reg_n_0_ ),
        .O(\processor/id_alu_x_src [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair52" *) 
  LUT5 #(
    .INIT(32'h0220A020)) 
    \alu_x_src[2]_i_1 
       (.I0(\processor/decode/instruction_reg_n_0_[5] ),
        .I1(\processor/decode/instruction_reg_n_0_[3] ),
        .I2(\processor/decode/instruction_reg_n_0_[6] ),
        .I3(\processor/decode/instruction_reg_n_0_ ),
        .I4(\processor/decode/instruction_reg_n_0_[4] ),
        .O(\processor/id_alu_x_src [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1A1A101023230111)) 
    \alu_y_src[0]_i_1 
       (.I0(\processor/decode/instruction_reg_n_0_[6] ),
        .I1(\processor/decode/instruction_reg_n_0_[3] ),
        .I2(\processor/decode/instruction_reg_n_0_[4] ),
        .I3(alu_y_src),
        .I4(\processor/decode/instruction_reg_n_0_[5] ),
        .I5(\processor/decode/instruction_reg_n_0_ ),
        .O(\processor/id_alu_y_src [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \alu_y_src[0]_i_2 
       (.I0(\processor/id_funct3 [0]),
        .I1(\processor/id_funct3 [1]),
        .O(alu_y_src));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \alu_y_src[1]_i_1 
       (.I0(\immediate[30]_i_2_n_0 ),
        .I1(\processor/id_funct3 [1]),
        .I2(\processor/id_funct3 [0]),
        .I3(\processor/decode/instruction_reg_n_0_[4] ),
        .I4(\processor/decode/instruction_reg_n_0_[5] ),
        .I5(\processor/decode/instruction_reg_n_0_ ),
        .O(\processor/id_alu_y_src [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00088808)) 
    \alu_y_src[2]_i_1 
       (.I0(\processor/decode/instruction_reg_n_0_[6] ),
        .I1(\processor/decode/instruction_reg_n_0_[5] ),
        .I2(\processor/decode/instruction_reg_n_0_[3] ),
        .I3(\processor/decode/instruction_reg_n_0_ ),
        .I4(\processor/decode/instruction_reg_n_0_[4] ),
        .O(\processor/id_alu_y_src [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \arbiter/FSM_sequential_state_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(FSM_sequential_state),
        .Q(\arbiter/state [0]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \arbiter/FSM_sequential_state_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\FSM_sequential_state[1]_i_1_n_0 ),
        .Q(\arbiter/state [1]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \arbiter/m1_inputs[ack] 
       (.I0(\arbiter/state [1]),
        .I1(\arbiter/state [0]),
        .I2(wb_ack_in),
        .O(icache_inputs));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \arbiter/m2_inputs[ack] 
       (.I0(\arbiter/state [0]),
        .I1(wb_ack_in),
        .I2(\arbiter/state [1]),
        .O(dmem_if_inputs));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[10]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [10]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [10]),
        .O(wb_adr_out[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[11]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [11]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [11]),
        .O(wb_adr_out[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[12]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [12]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [12]),
        .O(wb_adr_out[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[13]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [13]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [13]),
        .O(wb_adr_out[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[14]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [14]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [14]),
        .O(wb_adr_out[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[15]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [15]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [15]),
        .O(wb_adr_out[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[16]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [16]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [16]),
        .O(wb_adr_out[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[17]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [17]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [17]),
        .O(wb_adr_out[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[18]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [18]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [18]),
        .O(wb_adr_out[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[19]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [19]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [19]),
        .O(wb_adr_out[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[20]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [20]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [20]),
        .O(wb_adr_out[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[21]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [21]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [21]),
        .O(wb_adr_out[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[22]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [22]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [22]),
        .O(wb_adr_out[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[23]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [23]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [23]),
        .O(wb_adr_out[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[24]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [24]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [24]),
        .O(wb_adr_out[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[25]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [25]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [25]),
        .O(wb_adr_out[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[26]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [26]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [26]),
        .O(wb_adr_out[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[27]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [27]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [27]),
        .O(wb_adr_out[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[28]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [28]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [28]),
        .O(wb_adr_out[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[29]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [29]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [29]),
        .O(wb_adr_out[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[2]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [2]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [2]),
        .O(wb_adr_out[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[30]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [30]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [30]),
        .O(wb_adr_out[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[31]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [31]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [31]),
        .O(wb_adr_out[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[3]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [3]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [3]),
        .O(wb_adr_out[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[4]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [4]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [4]),
        .O(wb_adr_out[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[5]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [5]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [5]),
        .O(wb_adr_out[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[6]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [6]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [6]),
        .O(wb_adr_out[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[7]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [7]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [7]),
        .O(wb_adr_out[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[8]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [8]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [8]),
        .O(wb_adr_out[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_adr_out[9]_INST_0 
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[adr] [9]),
        .I2(\arbiter/state [0]),
        .I3(\icache_outputs[adr] [9]),
        .O(wb_adr_out[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_cyc_out 
       (.I0(icache_outputs),
        .I1(\arbiter/state [0]),
        .I2(dmem_if_outputs),
        .I3(\arbiter/state [1]),
        .O(wb_cyc_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_sel_out[0]_INST_0 
       (.I0(\icache_outputs[sel] ),
        .I1(\arbiter/state [0]),
        .I2(\dmem_if_outputs[sel] [0]),
        .I3(\arbiter/state [1]),
        .O(wb_sel_out[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_sel_out[1]_INST_0 
       (.I0(\icache_outputs[sel] ),
        .I1(\arbiter/state [0]),
        .I2(\dmem_if_outputs[sel] [1]),
        .I3(\arbiter/state [1]),
        .O(wb_sel_out[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_sel_out[2]_INST_0 
       (.I0(\icache_outputs[sel] ),
        .I1(\arbiter/state [0]),
        .I2(\dmem_if_outputs[sel] [2]),
        .I3(\arbiter/state [1]),
        .O(wb_sel_out[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_sel_out[3]_INST_0 
       (.I0(\icache_outputs[sel] ),
        .I1(\arbiter/state [0]),
        .I2(\dmem_if_outputs[sel] [3]),
        .I3(\arbiter/state [1]),
        .O(wb_sel_out[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \arbiter/wb_stb_out 
       (.I0(\icache_outputs[stb] ),
        .I1(\arbiter/state [0]),
        .I2(dmem_if_outputs),
        .I3(\arbiter/state [1]),
        .O(wb_stb_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h20000020)) 
    \branch[0]_i_1 
       (.I0(\processor/decode/instruction_reg_n_0_[5] ),
        .I1(\processor/decode/instruction_reg_n_0_[4] ),
        .I2(\processor/decode/instruction_reg_n_0_[6] ),
        .I3(\processor/decode/instruction_reg_n_0_ ),
        .I4(\processor/decode/instruction_reg_n_0_[3] ),
        .O(\processor/id_branch [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h1000)) 
    \branch[1]_i_1 
       (.I0(\processor/decode/instruction_reg_n_0_[3] ),
        .I1(\processor/decode/instruction_reg_n_0_[4] ),
        .I2(\processor/decode/instruction_reg_n_0_[6] ),
        .I3(\processor/decode/instruction_reg_n_0_[5] ),
        .O(\processor/id_branch [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \branch[2]_i_1 
       (.I0(\processor/id_shamt [1]),
        .I1(\processor/decode/instruction_reg_n_0_[3] ),
        .I2(\processor/id_shamt [3]),
        .I3(\processor/id_shamt [0]),
        .I4(branch),
        .I5(\branch[2]_i_3_n_0 ),
        .O(\processor/id_branch [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBFFFFFFF)) 
    \branch[2]_i_2 
       (.I0(\branch[2]_i_4_n_0 ),
        .I1(\processor/decode/instruction_reg_n_0_[4] ),
        .I2(\processor/decode/instruction_reg_n_0_[6] ),
        .I3(\processor/decode/instruction_reg_n_0_[5] ),
        .I4(data0[28]),
        .O(branch));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \branch[2]_i_3 
       (.I0(rd_write_out_i_2_n_0),
        .I1(data0[29]),
        .I2(\processor/id_shamt [2]),
        .I3(data0[31]),
        .I4(data0[30]),
        .O(\branch[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \branch[2]_i_4 
       (.I0(data0[26]),
        .I1(data0[27]),
        .I2(\processor/id_shamt [4]),
        .I3(data0[25]),
        .O(\branch[2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE200)) 
    cache_hit_i_1
       (.I0(cache_hit_i_2_n_0),
        .I1(imem_address[10]),
        .I2(cache_hit_i_3_n_0),
        .I3(\icache/to_std_logic ),
        .O(\icache/cache_hit0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_2
       (.I0(cache_hit_reg_i_4_n_0),
        .I1(cache_hit_reg_i_5_n_0),
        .I2(imem_address[9]),
        .I3(cache_hit_reg_i_6_n_0),
        .I4(imem_address[8]),
        .I5(cache_hit_reg_i_7_n_0),
        .O(cache_hit_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_28
       (.I0(\icache/valid [51]),
        .I1(\icache/valid [50]),
        .I2(imem_address[5]),
        .I3(\icache/valid [49]),
        .I4(imem_address[4]),
        .I5(\icache/valid [48]),
        .O(cache_hit_i_28_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_29
       (.I0(\icache/valid [55]),
        .I1(\icache/valid [54]),
        .I2(imem_address[5]),
        .I3(\icache/valid [53]),
        .I4(imem_address[4]),
        .I5(\icache/valid [52]),
        .O(cache_hit_i_29_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_3
       (.I0(cache_hit_reg_i_8_n_0),
        .I1(cache_hit_reg_i_9_n_0),
        .I2(imem_address[9]),
        .I3(cache_hit_reg_i_10_n_0),
        .I4(imem_address[8]),
        .I5(cache_hit_reg_i_11_n_0),
        .O(cache_hit_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_30
       (.I0(\icache/valid [59]),
        .I1(\icache/valid [58]),
        .I2(imem_address[5]),
        .I3(\icache/valid [57]),
        .I4(imem_address[4]),
        .I5(\icache/valid [56]),
        .O(cache_hit_i_30_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_31
       (.I0(\icache/valid [63]),
        .I1(\icache/valid [62]),
        .I2(imem_address[5]),
        .I3(\icache/valid [61]),
        .I4(imem_address[4]),
        .I5(\icache/valid [60]),
        .O(cache_hit_i_31_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_32
       (.I0(\icache/valid [35]),
        .I1(\icache/valid [34]),
        .I2(imem_address[5]),
        .I3(\icache/valid [33]),
        .I4(imem_address[4]),
        .I5(\icache/valid [32]),
        .O(cache_hit_i_32_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_33
       (.I0(\icache/valid [39]),
        .I1(\icache/valid [38]),
        .I2(imem_address[5]),
        .I3(\icache/valid [37]),
        .I4(imem_address[4]),
        .I5(\icache/valid [36]),
        .O(cache_hit_i_33_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_34
       (.I0(\icache/valid [43]),
        .I1(\icache/valid [42]),
        .I2(imem_address[5]),
        .I3(\icache/valid [41]),
        .I4(imem_address[4]),
        .I5(\icache/valid [40]),
        .O(cache_hit_i_34_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_35
       (.I0(\icache/valid [47]),
        .I1(\icache/valid [46]),
        .I2(imem_address[5]),
        .I3(\icache/valid [45]),
        .I4(imem_address[4]),
        .I5(\icache/valid [44]),
        .O(cache_hit_i_35_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_36
       (.I0(\icache/valid [19]),
        .I1(\icache/valid [18]),
        .I2(imem_address[5]),
        .I3(\icache/valid [17]),
        .I4(imem_address[4]),
        .I5(\icache/valid [16]),
        .O(cache_hit_i_36_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_37
       (.I0(\icache/valid [23]),
        .I1(\icache/valid [22]),
        .I2(imem_address[5]),
        .I3(\icache/valid [21]),
        .I4(imem_address[4]),
        .I5(\icache/valid [20]),
        .O(cache_hit_i_37_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_38
       (.I0(\icache/valid [27]),
        .I1(\icache/valid [26]),
        .I2(imem_address[5]),
        .I3(\icache/valid [25]),
        .I4(imem_address[4]),
        .I5(\icache/valid [24]),
        .O(cache_hit_i_38_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_39
       (.I0(\icache/valid [31]),
        .I1(\icache/valid [30]),
        .I2(imem_address[5]),
        .I3(\icache/valid [29]),
        .I4(imem_address[4]),
        .I5(\icache/valid [28]),
        .O(cache_hit_i_39_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_40
       (.I0(\icache/valid [3]),
        .I1(\icache/valid [2]),
        .I2(imem_address[5]),
        .I3(\icache/valid [1]),
        .I4(imem_address[4]),
        .I5(\icache/valid [0]),
        .O(cache_hit_i_40_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_41
       (.I0(\icache/valid [7]),
        .I1(\icache/valid [6]),
        .I2(imem_address[5]),
        .I3(\icache/valid [5]),
        .I4(imem_address[4]),
        .I5(\icache/valid [4]),
        .O(cache_hit_i_41_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_42
       (.I0(\icache/valid [11]),
        .I1(\icache/valid [10]),
        .I2(imem_address[5]),
        .I3(\icache/valid [9]),
        .I4(imem_address[4]),
        .I5(\icache/valid [8]),
        .O(cache_hit_i_42_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_43
       (.I0(\icache/valid [15]),
        .I1(\icache/valid [14]),
        .I2(imem_address[5]),
        .I3(\icache/valid [13]),
        .I4(imem_address[4]),
        .I5(\icache/valid [12]),
        .O(cache_hit_i_43_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_44
       (.I0(\icache/valid [115]),
        .I1(\icache/valid [114]),
        .I2(imem_address[5]),
        .I3(\icache/valid [113]),
        .I4(imem_address[4]),
        .I5(\icache/valid [112]),
        .O(cache_hit_i_44_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_45
       (.I0(\icache/valid [119]),
        .I1(\icache/valid [118]),
        .I2(imem_address[5]),
        .I3(\icache/valid [117]),
        .I4(imem_address[4]),
        .I5(\icache/valid [116]),
        .O(cache_hit_i_45_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_46
       (.I0(\icache/valid [123]),
        .I1(\icache/valid [122]),
        .I2(imem_address[5]),
        .I3(\icache/valid [121]),
        .I4(imem_address[4]),
        .I5(\icache/valid [120]),
        .O(cache_hit_i_46_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_47
       (.I0(\icache/valid [127]),
        .I1(\icache/valid [126]),
        .I2(imem_address[5]),
        .I3(\icache/valid [125]),
        .I4(imem_address[4]),
        .I5(\icache/valid [124]),
        .O(cache_hit_i_47_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_48
       (.I0(\icache/valid [99]),
        .I1(\icache/valid [98]),
        .I2(imem_address[5]),
        .I3(\icache/valid [97]),
        .I4(imem_address[4]),
        .I5(\icache/valid [96]),
        .O(cache_hit_i_48_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_49
       (.I0(\icache/valid [103]),
        .I1(\icache/valid [102]),
        .I2(imem_address[5]),
        .I3(\icache/valid [101]),
        .I4(imem_address[4]),
        .I5(\icache/valid [100]),
        .O(cache_hit_i_49_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_50
       (.I0(\icache/valid [107]),
        .I1(\icache/valid [106]),
        .I2(imem_address[5]),
        .I3(\icache/valid [105]),
        .I4(imem_address[4]),
        .I5(\icache/valid [104]),
        .O(cache_hit_i_50_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_51
       (.I0(\icache/valid [111]),
        .I1(\icache/valid [110]),
        .I2(imem_address[5]),
        .I3(\icache/valid [109]),
        .I4(imem_address[4]),
        .I5(\icache/valid [108]),
        .O(cache_hit_i_51_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_52
       (.I0(\icache/valid [83]),
        .I1(\icache/valid [82]),
        .I2(imem_address[5]),
        .I3(\icache/valid [81]),
        .I4(imem_address[4]),
        .I5(\icache/valid [80]),
        .O(cache_hit_i_52_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_53
       (.I0(\icache/valid [87]),
        .I1(\icache/valid [86]),
        .I2(imem_address[5]),
        .I3(\icache/valid [85]),
        .I4(imem_address[4]),
        .I5(\icache/valid [84]),
        .O(cache_hit_i_53_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_54
       (.I0(\icache/valid [91]),
        .I1(\icache/valid [90]),
        .I2(imem_address[5]),
        .I3(\icache/valid [89]),
        .I4(imem_address[4]),
        .I5(\icache/valid [88]),
        .O(cache_hit_i_54_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_55
       (.I0(\icache/valid [95]),
        .I1(\icache/valid [94]),
        .I2(imem_address[5]),
        .I3(\icache/valid [93]),
        .I4(imem_address[4]),
        .I5(\icache/valid [92]),
        .O(cache_hit_i_55_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_56
       (.I0(\icache/valid [67]),
        .I1(\icache/valid [66]),
        .I2(imem_address[5]),
        .I3(\icache/valid [65]),
        .I4(imem_address[4]),
        .I5(\icache/valid [64]),
        .O(cache_hit_i_56_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_57
       (.I0(\icache/valid [71]),
        .I1(\icache/valid [70]),
        .I2(imem_address[5]),
        .I3(\icache/valid [69]),
        .I4(imem_address[4]),
        .I5(\icache/valid [68]),
        .O(cache_hit_i_57_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_58
       (.I0(\icache/valid [75]),
        .I1(\icache/valid [74]),
        .I2(imem_address[5]),
        .I3(\icache/valid [73]),
        .I4(imem_address[4]),
        .I5(\icache/valid [72]),
        .O(cache_hit_i_58_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    cache_hit_i_59
       (.I0(\icache/valid [79]),
        .I1(\icache/valid [78]),
        .I2(imem_address[5]),
        .I3(\icache/valid [77]),
        .I4(imem_address[4]),
        .I5(\icache/valid [76]),
        .O(cache_hit_i_59_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 cache_hit_reg_i_10
       (.I0(cache_hit_reg_i_24_n_0),
        .I1(cache_hit_reg_i_25_n_0),
        .O(cache_hit_reg_i_10_n_0),
        .S(imem_address[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 cache_hit_reg_i_11
       (.I0(cache_hit_reg_i_26_n_0),
        .I1(cache_hit_reg_i_27_n_0),
        .O(cache_hit_reg_i_11_n_0),
        .S(imem_address[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 cache_hit_reg_i_12
       (.I0(cache_hit_i_28_n_0),
        .I1(cache_hit_i_29_n_0),
        .O(cache_hit_reg_i_12_n_0),
        .S(imem_address[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 cache_hit_reg_i_13
       (.I0(cache_hit_i_30_n_0),
        .I1(cache_hit_i_31_n_0),
        .O(cache_hit_reg_i_13_n_0),
        .S(imem_address[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 cache_hit_reg_i_14
       (.I0(cache_hit_i_32_n_0),
        .I1(cache_hit_i_33_n_0),
        .O(cache_hit_reg_i_14_n_0),
        .S(imem_address[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 cache_hit_reg_i_15
       (.I0(cache_hit_i_34_n_0),
        .I1(cache_hit_i_35_n_0),
        .O(cache_hit_reg_i_15_n_0),
        .S(imem_address[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 cache_hit_reg_i_16
       (.I0(cache_hit_i_36_n_0),
        .I1(cache_hit_i_37_n_0),
        .O(cache_hit_reg_i_16_n_0),
        .S(imem_address[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 cache_hit_reg_i_17
       (.I0(cache_hit_i_38_n_0),
        .I1(cache_hit_i_39_n_0),
        .O(cache_hit_reg_i_17_n_0),
        .S(imem_address[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 cache_hit_reg_i_18
       (.I0(cache_hit_i_40_n_0),
        .I1(cache_hit_i_41_n_0),
        .O(cache_hit_reg_i_18_n_0),
        .S(imem_address[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 cache_hit_reg_i_19
       (.I0(cache_hit_i_42_n_0),
        .I1(cache_hit_i_43_n_0),
        .O(cache_hit_reg_i_19_n_0),
        .S(imem_address[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 cache_hit_reg_i_20
       (.I0(cache_hit_i_44_n_0),
        .I1(cache_hit_i_45_n_0),
        .O(cache_hit_reg_i_20_n_0),
        .S(imem_address[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 cache_hit_reg_i_21
       (.I0(cache_hit_i_46_n_0),
        .I1(cache_hit_i_47_n_0),
        .O(cache_hit_reg_i_21_n_0),
        .S(imem_address[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 cache_hit_reg_i_22
       (.I0(cache_hit_i_48_n_0),
        .I1(cache_hit_i_49_n_0),
        .O(cache_hit_reg_i_22_n_0),
        .S(imem_address[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 cache_hit_reg_i_23
       (.I0(cache_hit_i_50_n_0),
        .I1(cache_hit_i_51_n_0),
        .O(cache_hit_reg_i_23_n_0),
        .S(imem_address[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 cache_hit_reg_i_24
       (.I0(cache_hit_i_52_n_0),
        .I1(cache_hit_i_53_n_0),
        .O(cache_hit_reg_i_24_n_0),
        .S(imem_address[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 cache_hit_reg_i_25
       (.I0(cache_hit_i_54_n_0),
        .I1(cache_hit_i_55_n_0),
        .O(cache_hit_reg_i_25_n_0),
        .S(imem_address[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 cache_hit_reg_i_26
       (.I0(cache_hit_i_56_n_0),
        .I1(cache_hit_i_57_n_0),
        .O(cache_hit_reg_i_26_n_0),
        .S(imem_address[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 cache_hit_reg_i_27
       (.I0(cache_hit_i_58_n_0),
        .I1(cache_hit_i_59_n_0),
        .O(cache_hit_reg_i_27_n_0),
        .S(imem_address[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 cache_hit_reg_i_4
       (.I0(cache_hit_reg_i_12_n_0),
        .I1(cache_hit_reg_i_13_n_0),
        .O(cache_hit_reg_i_4_n_0),
        .S(imem_address[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 cache_hit_reg_i_5
       (.I0(cache_hit_reg_i_14_n_0),
        .I1(cache_hit_reg_i_15_n_0),
        .O(cache_hit_reg_i_5_n_0),
        .S(imem_address[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 cache_hit_reg_i_6
       (.I0(cache_hit_reg_i_16_n_0),
        .I1(cache_hit_reg_i_17_n_0),
        .O(cache_hit_reg_i_6_n_0),
        .S(imem_address[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 cache_hit_reg_i_7
       (.I0(cache_hit_reg_i_18_n_0),
        .I1(cache_hit_reg_i_19_n_0),
        .O(cache_hit_reg_i_7_n_0),
        .S(imem_address[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 cache_hit_reg_i_8
       (.I0(cache_hit_reg_i_20_n_0),
        .I1(cache_hit_reg_i_21_n_0),
        .O(cache_hit_reg_i_8_n_0),
        .S(imem_address[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 cache_hit_reg_i_9
       (.I0(cache_hit_reg_i_22_n_0),
        .I1(cache_hit_reg_i_23_n_0),
        .O(cache_hit_reg_i_9_n_0),
        .S(imem_address[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    cache_memory_reg_0_i_1
       (.I0(pc[10]),
        .I1(pc_next[10]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0F0E)) 
    cancel_fetch_i_1
       (.I0(\mem_op[2]_i_5_n_0 ),
        .I1(\mem_op[2]_i_4_n_0 ),
        .I2(imem_ack),
        .I3(\processor/fetch/cancel_fetch ),
        .O(cancel_fetch_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h38)) 
    \cl_current_word[0]_i_1 
       (.I0(\icache/state_reg_n_0_[2] ),
        .I1(\cl_current_word[2]_i_2_n_0 ),
        .I2(\icache/cl_current_word_reg_n_0_ ),
        .O(cl_current_word));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair10" *) 
  LUT4 #(
    .INIT(16'h2F80)) 
    \cl_current_word[1]_i_1 
       (.I0(\icache/state_reg_n_0_[2] ),
        .I1(\icache/cl_current_word_reg_n_0_ ),
        .I2(\cl_current_word[2]_i_2_n_0 ),
        .I3(\icache/cl_current_word_reg_n_0_[1] ),
        .O(\cl_current_word[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair10" *) 
  LUT5 #(
    .INIT(32'h2AFF8000)) 
    \cl_current_word[2]_i_1 
       (.I0(\icache/state_reg_n_0_[2] ),
        .I1(\icache/cl_current_word_reg_n_0_[1] ),
        .I2(\icache/cl_current_word_reg_n_0_ ),
        .I3(\cl_current_word[2]_i_2_n_0 ),
        .I4(\icache/cl_current_word_reg_n_0_[2] ),
        .O(\cl_current_word[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000CC010001)) 
    \cl_current_word[2]_i_2 
       (.I0(\icache/cache_hit ),
        .I1(\icache/state_reg_n_0_[2] ),
        .I2(\icache/state_reg_n_0_[1] ),
        .I3(\icache/state_reg_n_0_ ),
        .I4(\cl_current_word[2]_i_3_n_0 ),
        .I5(reset),
        .O(\cl_current_word[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0808080800080808)) 
    \cl_current_word[2]_i_3 
       (.I0(wb_ack_in),
        .I1(\arbiter/state [0]),
        .I2(\arbiter/state [1]),
        .I3(\icache/cl_current_word_reg_n_0_[1] ),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .I5(\icache/cl_current_word_reg_n_0_[2] ),
        .O(\cl_current_word[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \cl_load_address[11]_i_1 
       (.I0(pc[11]),
        .I1(pc_next[11]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair138" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \cl_load_address[12]_i_1 
       (.I0(pc[12]),
        .I1(pc_next[12]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \cl_load_address[13]_i_1 
       (.I0(\icache/state_reg_n_0_[1] ),
        .I1(\icache/cache_hit ),
        .I2(\icache/state_reg_n_0_[2] ),
        .I3(\icache/state_reg_n_0_ ),
        .I4(reset),
        .O(cl_load_address));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair138" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \cl_load_address[13]_i_2 
       (.I0(pc[13]),
        .I1(pc_next[13]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \cl_load_address[14]_i_1 
       (.I0(pc[14]),
        .I1(pc_next[14]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \cl_load_address[15]_i_1 
       (.I0(pc[15]),
        .I1(pc_next[15]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \cl_load_address[16]_i_1 
       (.I0(pc[16]),
        .I1(pc_next[16]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \cl_load_address[17]_i_1 
       (.I0(pc[17]),
        .I1(pc_next[17]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair133" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \cl_load_address[18]_i_1 
       (.I0(pc[18]),
        .I1(pc_next[18]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair133" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \cl_load_address[19]_i_1 
       (.I0(pc[19]),
        .I1(pc_next[19]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \cl_load_address[20]_i_1 
       (.I0(pc[20]),
        .I1(pc_next[20]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \cl_load_address[21]_i_1 
       (.I0(pc[21]),
        .I1(pc_next[21]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \cl_load_address[22]_i_1 
       (.I0(pc[22]),
        .I1(pc_next[22]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \cl_load_address[23]_i_1 
       (.I0(pc[23]),
        .I1(pc_next[23]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair99" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \cl_load_address[24]_i_1 
       (.I0(pc[24]),
        .I1(pc_next[24]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair99" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \cl_load_address[25]_i_1 
       (.I0(pc[25]),
        .I1(pc_next[25]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \cl_load_address[26]_i_1 
       (.I0(pc[26]),
        .I1(pc_next[26]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \cl_load_address[27]_i_1 
       (.I0(pc[27]),
        .I1(pc_next[27]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair91" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \cl_load_address[28]_i_1 
       (.I0(pc[28]),
        .I1(pc_next[28]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \cl_load_address[29]_i_1 
       (.I0(pc[29]),
        .I1(pc_next[29]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \cl_load_address[30]_i_1 
       (.I0(pc[30]),
        .I1(pc_next[30]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair91" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \cl_load_address[31]_i_1 
       (.I0(pc[31]),
        .I1(pc_next[31]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    count_instr_out_i_1
       (.I0(reset),
        .I1(\processor/memory/p_1_in ),
        .I2(\mem_op[2]_i_5_n_0 ),
        .O(count_instr_out_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    count_instruction_i_1
       (.I0(imem_ack),
        .I1(\processor/execute/exception_taken0 ),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\mem_op[2]_i_5_n_0 ),
        .I4(\mem_op[2]_i_4_n_0 ),
        .I5(reset),
        .O(count_instruction_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \counter_mtime[0]_i_5 
       (.I0(\processor/csr_unit/counter_mtime_reg [0]),
        .O(counter_mtime));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \counter_mtime_reg[0]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO(counter_mtime_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .O({\counter_mtime_reg[0]_i_1_n_4 ,\counter_mtime_reg[0]_i_1_n_5 ,\counter_mtime_reg[0]_i_1_n_6 ,\counter_mtime_reg[0]_i_1_n_7 }),
        .S({\processor/csr_unit/counter_mtime_reg [3:1],counter_mtime}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \counter_mtime_reg[12]_i_1 
       (.CI(\counter_mtime_reg[8]_i_1_n_0 ),
        .CO({\counter_mtime_reg[12]_i_1_n_0 ,\counter_mtime_reg[12]_i_1_n_1 ,\counter_mtime_reg[12]_i_1_n_2 ,\counter_mtime_reg[12]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\counter_mtime_reg[12]_i_1_n_4 ,\counter_mtime_reg[12]_i_1_n_5 ,\counter_mtime_reg[12]_i_1_n_6 ,\counter_mtime_reg[12]_i_1_n_7 }),
        .S(\processor/csr_unit/counter_mtime_reg [15:12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \counter_mtime_reg[16]_i_1 
       (.CI(\counter_mtime_reg[12]_i_1_n_0 ),
        .CO({\counter_mtime_reg[16]_i_1_n_0 ,\counter_mtime_reg[16]_i_1_n_1 ,\counter_mtime_reg[16]_i_1_n_2 ,\counter_mtime_reg[16]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\counter_mtime_reg[16]_i_1_n_4 ,\counter_mtime_reg[16]_i_1_n_5 ,\counter_mtime_reg[16]_i_1_n_6 ,\counter_mtime_reg[16]_i_1_n_7 }),
        .S(\processor/csr_unit/counter_mtime_reg [19:16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \counter_mtime_reg[20]_i_1 
       (.CI(\counter_mtime_reg[16]_i_1_n_0 ),
        .CO({\counter_mtime_reg[20]_i_1_n_0 ,\counter_mtime_reg[20]_i_1_n_1 ,\counter_mtime_reg[20]_i_1_n_2 ,\counter_mtime_reg[20]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\counter_mtime_reg[20]_i_1_n_4 ,\counter_mtime_reg[20]_i_1_n_5 ,\counter_mtime_reg[20]_i_1_n_6 ,\counter_mtime_reg[20]_i_1_n_7 }),
        .S(\processor/csr_unit/counter_mtime_reg [23:20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \counter_mtime_reg[24]_i_1 
       (.CI(\counter_mtime_reg[20]_i_1_n_0 ),
        .CO({\counter_mtime_reg[24]_i_1_n_0 ,\counter_mtime_reg[24]_i_1_n_1 ,\counter_mtime_reg[24]_i_1_n_2 ,\counter_mtime_reg[24]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\counter_mtime_reg[24]_i_1_n_4 ,\counter_mtime_reg[24]_i_1_n_5 ,\counter_mtime_reg[24]_i_1_n_6 ,\counter_mtime_reg[24]_i_1_n_7 }),
        .S(\processor/csr_unit/counter_mtime_reg [27:24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \counter_mtime_reg[28]_i_1 
       (.CI(\counter_mtime_reg[24]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\counter_mtime_reg[28]_i_1_n_4 ,\counter_mtime_reg[28]_i_1_n_5 ,\counter_mtime_reg[28]_i_1_n_6 ,\counter_mtime_reg[28]_i_1_n_7 }),
        .S(\processor/csr_unit/counter_mtime_reg [31:28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \counter_mtime_reg[4]_i_1 
       (.CI(counter_mtime_reg[3]),
        .CO({\counter_mtime_reg[4]_i_1_n_0 ,\counter_mtime_reg[4]_i_1_n_1 ,\counter_mtime_reg[4]_i_1_n_2 ,\counter_mtime_reg[4]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\counter_mtime_reg[4]_i_1_n_4 ,\counter_mtime_reg[4]_i_1_n_5 ,\counter_mtime_reg[4]_i_1_n_6 ,\counter_mtime_reg[4]_i_1_n_7 }),
        .S(\processor/csr_unit/counter_mtime_reg [7:4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \counter_mtime_reg[8]_i_1 
       (.CI(\counter_mtime_reg[4]_i_1_n_0 ),
        .CO({\counter_mtime_reg[8]_i_1_n_0 ,\counter_mtime_reg[8]_i_1_n_1 ,\counter_mtime_reg[8]_i_1_n_2 ,\counter_mtime_reg[8]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\counter_mtime_reg[8]_i_1_n_4 ,\counter_mtime_reg[8]_i_1_n_5 ,\counter_mtime_reg[8]_i_1_n_6 ,\counter_mtime_reg[8]_i_1_n_7 }),
        .S(\processor/csr_unit/counter_mtime_reg [11:8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \csr_addr[0]_i_1 
       (.I0(csr_read_address_p[0]),
        .I1(\processor/decode/csr_addr__40 [0]),
        .I2(\processor/execute/exception_taken0 ),
        .O(csr_addr));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hC000AAAA)) 
    \csr_addr[10]_i_1 
       (.I0(csr_read_address_p[10]),
        .I1(\csr_addr[10]_i_2_n_0 ),
        .I2(data0[30]),
        .I3(\csr_addr[11]_i_2_n_0 ),
        .I4(\processor/execute/exception_taken0 ),
        .O(\csr_addr[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h1001B101)) 
    \csr_addr[10]_i_2 
       (.I0(\processor/decode/instruction_reg_n_0_ ),
        .I1(\processor/decode/instruction_reg_n_0_[3] ),
        .I2(\processor/decode/instruction_reg_n_0_[6] ),
        .I3(\processor/decode/instruction_reg_n_0_[5] ),
        .I4(\processor/decode/instruction_reg_n_0_[4] ),
        .O(\csr_addr[10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hC0AA)) 
    \csr_addr[11]_i_1 
       (.I0(csr_read_address_p[11]),
        .I1(\processor/id_immediate [11]),
        .I2(\csr_addr[11]_i_2_n_0 ),
        .I3(\processor/execute/exception_taken0 ),
        .O(\csr_addr[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \csr_addr[11]_i_2 
       (.I0(\csr_addr[11]_i_3_n_0 ),
        .I1(\csr_read_address_p[0]_i_3_n_0 ),
        .I2(\processor/id_immediate [0]),
        .I3(\processor/id_immediate [1]),
        .I4(\csr_addr[11]_i_4_n_0 ),
        .O(\csr_addr[11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFDFFFF)) 
    \csr_addr[11]_i_3 
       (.I0(data0[28]),
        .I1(data0[30]),
        .I2(\processor/id_immediate [11]),
        .I3(data0[29]),
        .I4(\csr_addr[10]_i_2_n_0 ),
        .O(\csr_addr[11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFEF0F0)) 
    \csr_addr[11]_i_4 
       (.I0(data0[26]),
        .I1(data0[27]),
        .I2(\processor/id_immediate [4]),
        .I3(data0[25]),
        .I4(\csr_addr[10]_i_2_n_0 ),
        .O(\csr_addr[11]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hC0AA)) 
    \csr_addr[1]_i_1 
       (.I0(csr_read_address_p[1]),
        .I1(\processor/id_immediate [1]),
        .I2(\csr_addr[11]_i_2_n_0 ),
        .I3(\processor/execute/exception_taken0 ),
        .O(\csr_addr[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hC0AA)) 
    \csr_addr[2]_i_1 
       (.I0(csr_read_address_p[2]),
        .I1(\processor/id_immediate [2]),
        .I2(\csr_addr[11]_i_2_n_0 ),
        .I3(\processor/execute/exception_taken0 ),
        .O(\csr_addr[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hC0AA)) 
    \csr_addr[3]_i_1 
       (.I0(csr_read_address_p[3]),
        .I1(\processor/id_immediate [3]),
        .I2(\csr_addr[11]_i_2_n_0 ),
        .I3(\processor/execute/exception_taken0 ),
        .O(\csr_addr[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hC0AA)) 
    \csr_addr[4]_i_1 
       (.I0(csr_read_address_p[4]),
        .I1(\processor/id_immediate [4]),
        .I2(\csr_addr[11]_i_2_n_0 ),
        .I3(\processor/execute/exception_taken0 ),
        .O(\csr_addr[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hC000AAAA)) 
    \csr_addr[5]_i_1 
       (.I0(csr_read_address_p[5]),
        .I1(\csr_addr[10]_i_2_n_0 ),
        .I2(data0[25]),
        .I3(\csr_addr[11]_i_2_n_0 ),
        .I4(\processor/execute/exception_taken0 ),
        .O(\csr_addr[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF8F8FF00)) 
    \csr_addr[6]_i_1 
       (.I0(\csr_addr[10]_i_2_n_0 ),
        .I1(data0[26]),
        .I2(\csr_addr[9]_i_2_n_0 ),
        .I3(csr_read_address_p[6]),
        .I4(\processor/execute/exception_taken0 ),
        .O(\csr_addr[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hC000AAAA)) 
    \csr_addr[7]_i_1 
       (.I0(csr_read_address_p[7]),
        .I1(\csr_addr[10]_i_2_n_0 ),
        .I2(data0[27]),
        .I3(\csr_addr[11]_i_2_n_0 ),
        .I4(\processor/execute/exception_taken0 ),
        .O(\csr_addr[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF8F8FF00)) 
    \csr_addr[8]_i_1 
       (.I0(\csr_addr[10]_i_2_n_0 ),
        .I1(data0[28]),
        .I2(\csr_addr[9]_i_2_n_0 ),
        .I3(csr_read_address_p[8]),
        .I4(\processor/execute/exception_taken0 ),
        .O(\csr_addr[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF8F8FF00)) 
    \csr_addr[9]_i_1 
       (.I0(\csr_addr[10]_i_2_n_0 ),
        .I1(data0[29]),
        .I2(\csr_addr[9]_i_2_n_0 ),
        .I3(csr_read_address_p[9]),
        .I4(\processor/execute/exception_taken0 ),
        .O(\csr_addr[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \csr_addr[9]_i_2 
       (.I0(\csr_addr[9]_i_3_n_0 ),
        .I1(\csr_read_address_p[0]_i_3_n_0 ),
        .I2(data0[28]),
        .I3(\csr_addr[10]_i_2_n_0 ),
        .I4(\processor/id_immediate [1]),
        .I5(\csr_addr[11]_i_4_n_0 ),
        .O(\csr_addr[9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFEFAFA)) 
    \csr_addr[9]_i_3 
       (.I0(\processor/id_immediate [11]),
        .I1(data0[30]),
        .I2(\processor/id_immediate [0]),
        .I3(data0[29]),
        .I4(\csr_addr[10]_i_2_n_0 ),
        .O(\csr_addr[9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \csr_addr_out[11]_i_1 
       (.I0(\processor/memory/p_1_in ),
        .I1(\mem_op[2]_i_5_n_0 ),
        .I2(reset),
        .O(csr_addr_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[0]_i_1 
       (.I0(\processor/ex_pc [0]),
        .I1(\processor/execute/csr_alu_instance/b [0]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[0]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(csr_data_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \csr_data_out[0]_i_2 
       (.I0(\processor/execute/rs1_addr [0]),
        .I1(\processor/execute/rs1_forwarded [0]),
        .I2(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00FE)) 
    \csr_data_out[0]_i_3 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\csr_data_out[0]_i_5_n_0 ),
        .I2(\csr_data_out[0]_i_6_n_0 ),
        .I3(\csr_data_out[0]_i_7_n_0 ),
        .O(\csr_data_out[0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[0]_i_4 
       (.I0(\processor/mem_rd_data [0]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [0]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [0]),
        .O(\processor/execute/rs1_forwarded [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000474700FF)) 
    \csr_data_out[0]_i_5 
       (.I0(\processor/wb_csr_data [0]),
        .I1(\csr_data_out[30]_i_8_n_0 ),
        .I2(\processor/csr_read_data [0]),
        .I3(\processor/wb_exception_context[badaddr] [0]),
        .I4(\csr_data_out[31]_i_21_n_0 ),
        .I5(\csr_data_out[4]_i_9_n_0 ),
        .O(\csr_data_out[0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4E004E0000004E00)) 
    \csr_data_out[0]_i_6 
       (.I0(\csr_data_out[30]_i_5_n_0 ),
        .I1(\csr_data_out[0]_i_8_n_0 ),
        .I2(\processor/mem_csr_data [0]),
        .I3(\csr_data_out[4]_i_9_n_0 ),
        .I4(\processor/wb_exception_context[ie] ),
        .I5(\csr_data_out[3]_i_9_n_0 ),
        .O(\csr_data_out[0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF44F444F444F4)) 
    \csr_data_out[0]_i_7 
       (.I0(\csr_data_out[31]_i_24_n_0 ),
        .I1(\processor/mem_exception_context[cause] [0]),
        .I2(\processor/mem_exception_context[badaddr] [0]),
        .I3(\csr_data_out[31]_i_25_n_0 ),
        .I4(\processor/mem_exception_context[ie] ),
        .I5(\csr_data_out[4]_i_11_n_0 ),
        .O(\csr_data_out[0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFDFFFFFFFFFFFFFF)) 
    \csr_data_out[0]_i_8 
       (.I0(\processor/wb_exception ),
        .I1(\processor/ex_csr_address [0]),
        .I2(\csr_data_out[30]_i_10_n_0 ),
        .I3(\processor/ex_csr_address[6]_repN_1 ),
        .I4(\processor/ex_csr_address [1]),
        .I5(\processor/wb_exception_context[cause] [0]),
        .O(\csr_data_out[0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[10]_i_1 
       (.I0(\processor/ex_pc [10]),
        .I1(\processor/execute/csr_alu_instance/b [10]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[10]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[10]_i_2 
       (.I0(\processor/execute/rs1_forwarded [10]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000F2F2F2)) 
    \csr_data_out[10]_i_3 
       (.I0(\csr_data_out[10]_i_5_n_0 ),
        .I1(\csr_data_out[10]_i_6_n_0 ),
        .I2(\csr_data_out[31]_i_6_n_0 ),
        .I3(\processor/mem_exception_context[badaddr] [10]),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\csr_data_out[11]_i_7_n_0 ),
        .O(\csr_data_out[10]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[10]_i_4 
       (.I0(\processor/mem_rd_data [10]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [10]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [10]),
        .O(\processor/execute/rs1_forwarded [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAABABFFFFFBABF)) 
    \csr_data_out[10]_i_5 
       (.I0(\csr_data_out[4]_i_9_n_0 ),
        .I1(\processor/wb_csr_data [10]),
        .I2(\csr_data_out[30]_i_8_n_0 ),
        .I3(\processor/csr_read_data [10]),
        .I4(\csr_data_out[30]_i_9_n_0 ),
        .I5(\processor/wb_exception_context[badaddr] [10]),
        .O(\csr_data_out[10]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFFFFFFA8000000)) 
    \csr_data_out[10]_i_6 
       (.I0(\processor/mem_csr_data [10]),
        .I1(\processor/mem_csr_write [1]),
        .I2(\processor/mem_csr_write [0]),
        .I3(\processor/execute/csr_value_forwarded30_out ),
        .I4(\processor/execute/csr_writeable ),
        .I5(\csr_data_out[31]_i_19_n_0 ),
        .O(\csr_data_out[10]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[11]_i_1 
       (.I0(\processor/ex_pc [11]),
        .I1(\processor/execute/csr_alu_instance/b [11]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[11]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[11]_i_2 
       (.I0(\processor/execute/rs1_forwarded [11]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000F2F2F2)) 
    \csr_data_out[11]_i_3 
       (.I0(\csr_data_out[11]_i_5_n_0 ),
        .I1(\csr_data_out[11]_i_6_n_0 ),
        .I2(\csr_data_out[31]_i_6_n_0 ),
        .I3(\processor/mem_exception_context[badaddr] [11]),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\csr_data_out[11]_i_7_n_0 ),
        .O(\csr_data_out[11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[11]_i_4 
       (.I0(\processor/mem_rd_data [11]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [11]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [11]),
        .O(\processor/execute/rs1_forwarded [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAABABFFFFFBABF)) 
    \csr_data_out[11]_i_5 
       (.I0(\csr_data_out[4]_i_9_n_0 ),
        .I1(\processor/wb_csr_data [11]),
        .I2(\csr_data_out[30]_i_8_n_0 ),
        .I3(\processor/csr_read_data [11]),
        .I4(\csr_data_out[30]_i_9_n_0 ),
        .I5(\processor/wb_exception_context[badaddr] [11]),
        .O(\csr_data_out[11]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFFFFFFA8000000)) 
    \csr_data_out[11]_i_6 
       (.I0(\processor/mem_csr_data [11]),
        .I1(\processor/mem_csr_write [1]),
        .I2(\processor/mem_csr_write [0]),
        .I3(\processor/execute/csr_value_forwarded30_out ),
        .I4(\processor/execute/csr_writeable ),
        .I5(\csr_data_out[31]_i_19_n_0 ),
        .O(\csr_data_out[11]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \csr_data_out[11]_i_7 
       (.I0(\processor/mem_exception ),
        .I1(\csr_data_out[11]_i_8_n_0 ),
        .I2(\processor/ex_csr_address [11]),
        .I3(\processor/ex_csr_address [2]),
        .I4(\processor/ex_csr_address [5]),
        .I5(\csr_data_out[31]_i_15_n_0 ),
        .O(\csr_data_out[11]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \csr_data_out[11]_i_8 
       (.I0(\processor/ex_csr_address [6]),
        .I1(\processor/ex_csr_address [0]),
        .I2(\processor/ex_csr_address [1]),
        .O(\csr_data_out[11]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[12]_i_1 
       (.I0(\processor/ex_pc [12]),
        .I1(\processor/execute/csr_alu_instance/b [12]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[12]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[12]_i_2 
       (.I0(\processor/execute/rs1_forwarded [12]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FF07FF07FF07)) 
    \csr_data_out[12]_i_3 
       (.I0(\csr_data_out[30]_i_5_n_0_repN ),
        .I1(\processor/mem_csr_data [12]),
        .I2(\csr_data_out[12]_i_5_n_0 ),
        .I3(\csr_data_out[31]_i_6_n_0 ),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\processor/mem_exception_context[badaddr] [12]),
        .O(\csr_data_out[12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[12]_i_4 
       (.I0(\processor/mem_rd_data [12]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [12]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [12]),
        .O(\processor/execute/rs1_forwarded [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFD800D8)) 
    \csr_data_out[12]_i_5 
       (.I0(\csr_data_out[30]_i_8_n_0 ),
        .I1(\processor/wb_csr_data [12]),
        .I2(\processor/csr_read_data [12]),
        .I3(\csr_data_out[30]_i_9_n_0 ),
        .I4(\processor/wb_exception_context[badaddr] [12]),
        .I5(\csr_data_out[4]_i_9_n_0 ),
        .O(\csr_data_out[12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[13]_i_1 
       (.I0(\processor/ex_pc [13]),
        .I1(\processor/execute/csr_alu_instance/b [13]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[13]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[13]_i_2 
       (.I0(\processor/execute/rs1_forwarded [13]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FF07FF07FF07)) 
    \csr_data_out[13]_i_3 
       (.I0(\csr_data_out[30]_i_5_n_0 ),
        .I1(\processor/mem_csr_data [13]),
        .I2(\csr_data_out[13]_i_5_n_0 ),
        .I3(\csr_data_out[31]_i_6_n_0 ),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\processor/mem_exception_context[badaddr] [13]),
        .O(\csr_data_out[13]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[13]_i_4 
       (.I0(\processor/mem_rd_data [13]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [13]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [13]),
        .O(\processor/execute/rs1_forwarded [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFD800D8)) 
    \csr_data_out[13]_i_5 
       (.I0(\csr_data_out[30]_i_8_n_0 ),
        .I1(\processor/wb_csr_data [13]),
        .I2(\processor/csr_read_data [13]),
        .I3(\csr_data_out[30]_i_9_n_0 ),
        .I4(\processor/wb_exception_context[badaddr] [13]),
        .I5(\csr_data_out[4]_i_9_n_0 ),
        .O(\csr_data_out[13]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[14]_i_1 
       (.I0(\processor/ex_pc [14]),
        .I1(\processor/execute/csr_alu_instance/b [14]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[14]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[14]_i_2 
       (.I0(\processor/execute/rs1_forwarded [14]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FF07FF07FF07)) 
    \csr_data_out[14]_i_3 
       (.I0(\csr_data_out[30]_i_5_n_0_repN ),
        .I1(\processor/mem_csr_data [14]),
        .I2(\csr_data_out[14]_i_5_n_0 ),
        .I3(\csr_data_out[31]_i_6_n_0 ),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\processor/mem_exception_context[badaddr] [14]),
        .O(\csr_data_out[14]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[14]_i_4 
       (.I0(\processor/mem_rd_data [14]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [14]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [14]),
        .O(\processor/execute/rs1_forwarded [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFD800D8)) 
    \csr_data_out[14]_i_5 
       (.I0(\csr_data_out[30]_i_8_n_0 ),
        .I1(\processor/wb_csr_data [14]),
        .I2(\processor/csr_read_data [14]),
        .I3(\csr_data_out[30]_i_9_n_0 ),
        .I4(\processor/wb_exception_context[badaddr] [14]),
        .I5(\csr_data_out[4]_i_9_n_0 ),
        .O(\csr_data_out[14]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[15]_i_1 
       (.I0(\processor/ex_pc [15]),
        .I1(\processor/execute/csr_alu_instance/b [15]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[15]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[15]_i_2 
       (.I0(\processor/execute/rs1_forwarded [15]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FF07FF07FF07)) 
    \csr_data_out[15]_i_3 
       (.I0(\csr_data_out[30]_i_5_n_0 ),
        .I1(\processor/mem_csr_data [15]),
        .I2(\csr_data_out[15]_i_5_n_0 ),
        .I3(\csr_data_out[31]_i_6_n_0 ),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\processor/mem_exception_context[badaddr] [15]),
        .O(\csr_data_out[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[15]_i_4 
       (.I0(\processor/mem_rd_data [15]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [15]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [15]),
        .O(\processor/execute/rs1_forwarded [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFD800D8)) 
    \csr_data_out[15]_i_5 
       (.I0(\csr_data_out[30]_i_8_n_0 ),
        .I1(\processor/wb_csr_data [15]),
        .I2(\processor/csr_read_data [15]),
        .I3(\csr_data_out[30]_i_9_n_0 ),
        .I4(\processor/wb_exception_context[badaddr] [15]),
        .I5(\csr_data_out[4]_i_9_n_0 ),
        .O(\csr_data_out[15]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[16]_i_1 
       (.I0(\processor/ex_pc [16]),
        .I1(\processor/execute/csr_alu_instance/b [16]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[16]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[16]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[16]_i_2 
       (.I0(\processor/execute/rs1_forwarded [16]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FF07FF07FF07)) 
    \csr_data_out[16]_i_3 
       (.I0(\csr_data_out[30]_i_5_n_0 ),
        .I1(\processor/mem_csr_data [16]),
        .I2(\csr_data_out[16]_i_5_n_0 ),
        .I3(\csr_data_out[31]_i_6_n_0 ),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\processor/mem_exception_context[badaddr] [16]),
        .O(\csr_data_out[16]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[16]_i_4 
       (.I0(\processor/mem_rd_data [16]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [16]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [16]),
        .O(\processor/execute/rs1_forwarded [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFD800D8)) 
    \csr_data_out[16]_i_5 
       (.I0(\csr_data_out[30]_i_8_n_0 ),
        .I1(\processor/wb_csr_data [16]),
        .I2(\processor/csr_read_data [16]),
        .I3(\csr_data_out[30]_i_9_n_0 ),
        .I4(\processor/wb_exception_context[badaddr] [16]),
        .I5(\csr_data_out[4]_i_9_n_0 ),
        .O(\csr_data_out[16]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[17]_i_1 
       (.I0(\processor/ex_pc [17]),
        .I1(\processor/execute/csr_alu_instance/b [17]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[17]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[17]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[17]_i_2 
       (.I0(\processor/execute/rs1_forwarded [17]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FF07FF07FF07)) 
    \csr_data_out[17]_i_3 
       (.I0(\csr_data_out[30]_i_5_n_0 ),
        .I1(\processor/mem_csr_data [17]),
        .I2(\csr_data_out[17]_i_5_n_0 ),
        .I3(\csr_data_out[31]_i_6_n_0 ),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\processor/mem_exception_context[badaddr] [17]),
        .O(\csr_data_out[17]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[17]_i_4 
       (.I0(\processor/mem_rd_data [17]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [17]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [17]),
        .O(\processor/execute/rs1_forwarded [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFD800D8)) 
    \csr_data_out[17]_i_5 
       (.I0(\csr_data_out[30]_i_8_n_0 ),
        .I1(\processor/wb_csr_data [17]),
        .I2(\processor/csr_read_data [17]),
        .I3(\csr_data_out[30]_i_9_n_0 ),
        .I4(\processor/wb_exception_context[badaddr] [17]),
        .I5(\csr_data_out[4]_i_9_n_0 ),
        .O(\csr_data_out[17]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[18]_i_1 
       (.I0(\processor/ex_pc [18]),
        .I1(\processor/execute/csr_alu_instance/b [18]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[18]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[18]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[18]_i_2 
       (.I0(\processor/execute/rs1_forwarded [18]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FF07FF07FF07)) 
    \csr_data_out[18]_i_3 
       (.I0(\csr_data_out[30]_i_5_n_0 ),
        .I1(\processor/mem_csr_data [18]),
        .I2(\csr_data_out[18]_i_5_n_0 ),
        .I3(\csr_data_out[31]_i_6_n_0 ),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\processor/mem_exception_context[badaddr] [18]),
        .O(\csr_data_out[18]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[18]_i_4 
       (.I0(\processor/mem_rd_data [18]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [18]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [18]),
        .O(\processor/execute/rs1_forwarded [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFD800D8)) 
    \csr_data_out[18]_i_5 
       (.I0(\csr_data_out[30]_i_8_n_0 ),
        .I1(\processor/wb_csr_data [18]),
        .I2(\processor/csr_read_data [18]),
        .I3(\csr_data_out[30]_i_9_n_0 ),
        .I4(\processor/wb_exception_context[badaddr] [18]),
        .I5(\csr_data_out[4]_i_9_n_0 ),
        .O(\csr_data_out[18]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[19]_i_1 
       (.I0(\processor/ex_pc [19]),
        .I1(\processor/execute/csr_alu_instance/b [19]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[19]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[19]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[19]_i_2 
       (.I0(\processor/execute/rs1_forwarded [19]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FF07FF07FF07)) 
    \csr_data_out[19]_i_3 
       (.I0(\csr_data_out[30]_i_5_n_0 ),
        .I1(\processor/mem_csr_data [19]),
        .I2(\csr_data_out[19]_i_5_n_0 ),
        .I3(\csr_data_out[31]_i_6_n_0 ),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\processor/mem_exception_context[badaddr] [19]),
        .O(\csr_data_out[19]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[19]_i_4 
       (.I0(\processor/mem_rd_data [19]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [19]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [19]),
        .O(\processor/execute/rs1_forwarded [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFD800D8)) 
    \csr_data_out[19]_i_5 
       (.I0(\csr_data_out[30]_i_8_n_0 ),
        .I1(\processor/wb_csr_data [19]),
        .I2(\processor/csr_read_data [19]),
        .I3(\csr_data_out[30]_i_9_n_0 ),
        .I4(\processor/wb_exception_context[badaddr] [19]),
        .I5(\csr_data_out[4]_i_9_n_0 ),
        .O(\csr_data_out[19]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[1]_i_1 
       (.I0(\processor/ex_pc [1]),
        .I1(\processor/execute/csr_alu_instance/b [1]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[1]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \csr_data_out[1]_i_2 
       (.I0(\processor/execute/rs1_addr [1]),
        .I1(\processor/execute/rs1_forwarded [1]),
        .I2(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000EEEEEEFE)) 
    \csr_data_out[1]_i_3 
       (.I0(\csr_data_out[1]_i_5_n_0 ),
        .I1(\csr_data_out[31]_i_6_n_0 ),
        .I2(\csr_data_out[1]_i_6_n_0 ),
        .I3(\csr_data_out[1]_i_7_n_0 ),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\csr_data_out[1]_i_8_n_0 ),
        .O(\csr_data_out[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[1]_i_4 
       (.I0(\processor/mem_rd_data [1]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [1]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [1]),
        .O(\processor/execute/rs1_forwarded [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h110F111111111111)) 
    \csr_data_out[1]_i_5 
       (.I0(\csr_data_out[31]_i_16_n_0 ),
        .I1(\processor/wb_exception_context[cause] [1]),
        .I2(\processor/mem_csr_data [1]),
        .I3(\csr_data_out[31]_i_18_n_0 ),
        .I4(\processor/execute/csr_value_forwarded30_out ),
        .I5(\processor/execute/csr_writeable ),
        .O(\csr_data_out[1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1555D555FFFFFFFF)) 
    \csr_data_out[1]_i_6 
       (.I0(\processor/csr_read_data [1]),
        .I1(\processor/csr_unit/tohost_data1__0 ),
        .I2(\processor/execute/csr_value_forwarded3 ),
        .I3(\processor/execute/csr_writeable ),
        .I4(\processor/wb_csr_data [1]),
        .I5(\csr_data_out[31]_i_21_n_0 ),
        .O(\csr_data_out[1]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[1]_i_7 
       (.I0(\processor/wb_exception_context[badaddr] [1]),
        .I1(\csr_data_out[31]_i_21_n_0 ),
        .O(\csr_data_out[1]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \csr_data_out[1]_i_8 
       (.I0(\csr_data_out[31]_i_24_n_0 ),
        .I1(\processor/mem_exception_context[cause] [1]),
        .I2(\processor/mem_exception_context[badaddr] [1]),
        .I3(\csr_data_out[31]_i_25_n_0 ),
        .I4(\csr_data_out[4]_i_11_n_0 ),
        .O(\csr_data_out[1]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[20]_i_1 
       (.I0(\processor/ex_pc [20]),
        .I1(\processor/execute/csr_alu_instance/b [20]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[20]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[20]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[20]_i_2 
       (.I0(\processor/execute/rs1_forwarded [20]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FF07FF07FF07)) 
    \csr_data_out[20]_i_3 
       (.I0(\csr_data_out[30]_i_5_n_0 ),
        .I1(\processor/mem_csr_data [20]),
        .I2(\csr_data_out[20]_i_5_n_0 ),
        .I3(\csr_data_out[31]_i_6_n_0 ),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\processor/mem_exception_context[badaddr] [20]),
        .O(\csr_data_out[20]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[20]_i_4 
       (.I0(\processor/mem_rd_data [20]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [20]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [20]),
        .O(\processor/execute/rs1_forwarded [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFD800D8)) 
    \csr_data_out[20]_i_5 
       (.I0(\csr_data_out[30]_i_8_n_0 ),
        .I1(\processor/wb_csr_data [20]),
        .I2(\processor/csr_read_data [20]),
        .I3(\csr_data_out[30]_i_9_n_0 ),
        .I4(\processor/wb_exception_context[badaddr] [20]),
        .I5(\csr_data_out[4]_i_9_n_0 ),
        .O(\csr_data_out[20]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[21]_i_1 
       (.I0(\processor/ex_pc [21]),
        .I1(\processor/execute/csr_alu_instance/b [21]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[21]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[21]_i_2 
       (.I0(\processor/execute/rs1_forwarded [21]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FF07FF07FF07)) 
    \csr_data_out[21]_i_3 
       (.I0(\csr_data_out[30]_i_5_n_0 ),
        .I1(\processor/mem_csr_data [21]),
        .I2(\csr_data_out[21]_i_5_n_0 ),
        .I3(\csr_data_out[31]_i_6_n_0 ),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\processor/mem_exception_context[badaddr] [21]),
        .O(\csr_data_out[21]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[21]_i_4 
       (.I0(\processor/mem_rd_data [21]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [21]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [21]),
        .O(\processor/execute/rs1_forwarded [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFD800D8)) 
    \csr_data_out[21]_i_5 
       (.I0(\csr_data_out[30]_i_8_n_0 ),
        .I1(\processor/wb_csr_data [21]),
        .I2(\processor/csr_read_data [21]),
        .I3(\csr_data_out[30]_i_9_n_0 ),
        .I4(\processor/wb_exception_context[badaddr] [21]),
        .I5(\csr_data_out[4]_i_9_n_0 ),
        .O(\csr_data_out[21]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[22]_i_1 
       (.I0(\processor/ex_pc [22]),
        .I1(\processor/execute/csr_alu_instance/b [22]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[22]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[22]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[22]_i_2 
       (.I0(\processor/execute/rs1_forwarded [22]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FF07FF07FF07)) 
    \csr_data_out[22]_i_3 
       (.I0(\csr_data_out[30]_i_5_n_0 ),
        .I1(\processor/mem_csr_data [22]),
        .I2(\csr_data_out[22]_i_5_n_0 ),
        .I3(\csr_data_out[31]_i_6_n_0 ),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\processor/mem_exception_context[badaddr] [22]),
        .O(\csr_data_out[22]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[22]_i_4 
       (.I0(\processor/mem_rd_data [22]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [22]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [22]),
        .O(\processor/execute/rs1_forwarded [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFD800D8)) 
    \csr_data_out[22]_i_5 
       (.I0(\csr_data_out[30]_i_8_n_0 ),
        .I1(\processor/wb_csr_data [22]),
        .I2(\processor/csr_read_data [22]),
        .I3(\csr_data_out[30]_i_9_n_0 ),
        .I4(\processor/wb_exception_context[badaddr] [22]),
        .I5(\csr_data_out[4]_i_9_n_0 ),
        .O(\csr_data_out[22]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[23]_i_1 
       (.I0(\processor/ex_pc [23]),
        .I1(\processor/execute/csr_alu_instance/b [23]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[23]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[23]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[23]_i_2 
       (.I0(\processor/execute/rs1_forwarded [23]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FF07FF07FF07)) 
    \csr_data_out[23]_i_3 
       (.I0(\csr_data_out[30]_i_5_n_0 ),
        .I1(\processor/mem_csr_data [23]),
        .I2(\csr_data_out[23]_i_5_n_0 ),
        .I3(\csr_data_out[31]_i_6_n_0 ),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\processor/mem_exception_context[badaddr] [23]),
        .O(\csr_data_out[23]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[23]_i_4 
       (.I0(\processor/mem_rd_data [23]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [23]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [23]),
        .O(\processor/execute/rs1_forwarded [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFD800D8)) 
    \csr_data_out[23]_i_5 
       (.I0(\csr_data_out[30]_i_8_n_0 ),
        .I1(\processor/wb_csr_data [23]),
        .I2(\processor/csr_read_data [23]),
        .I3(\csr_data_out[30]_i_9_n_0 ),
        .I4(\processor/wb_exception_context[badaddr] [23]),
        .I5(\csr_data_out[4]_i_9_n_0 ),
        .O(\csr_data_out[23]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[24]_i_1 
       (.I0(\processor/ex_pc [24]),
        .I1(\processor/execute/csr_alu_instance/b [24]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[24]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[24]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[24]_i_2 
       (.I0(\processor/execute/rs1_forwarded [24]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FF07FF07FF07)) 
    \csr_data_out[24]_i_3 
       (.I0(\csr_data_out[30]_i_5_n_0 ),
        .I1(\processor/mem_csr_data [24]),
        .I2(\csr_data_out[24]_i_5_n_0 ),
        .I3(\csr_data_out[31]_i_6_n_0 ),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\processor/mem_exception_context[badaddr] [24]),
        .O(\csr_data_out[24]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[24]_i_4 
       (.I0(\processor/mem_rd_data [24]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [24]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [24]),
        .O(\processor/execute/rs1_forwarded [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    \csr_data_out[24]_i_5 
       (.I0(\processor/wb_csr_data [24]),
        .I1(\csr_data_out[30]_i_8_n_0 ),
        .I2(\processor/csr_read_data [24]),
        .I3(\csr_data_out[30]_i_9_n_0 ),
        .I4(\processor/wb_exception_context[badaddr] [24]),
        .I5(\csr_data_out[4]_i_9_n_0 ),
        .O(\csr_data_out[24]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[25]_i_1 
       (.I0(\processor/ex_pc [25]),
        .I1(\processor/execute/csr_alu_instance/b [25]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[25]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[25]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[25]_i_2 
       (.I0(\processor/execute/rs1_forwarded [25]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FF07FF07FF07)) 
    \csr_data_out[25]_i_3 
       (.I0(\csr_data_out[30]_i_5_n_0 ),
        .I1(\processor/mem_csr_data [25]),
        .I2(\csr_data_out[25]_i_5_n_0 ),
        .I3(\csr_data_out[31]_i_6_n_0 ),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\processor/mem_exception_context[badaddr] [25]),
        .O(\csr_data_out[25]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[25]_i_4 
       (.I0(\processor/mem_rd_data [25]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [25]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [25]),
        .O(\processor/execute/rs1_forwarded [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    \csr_data_out[25]_i_5 
       (.I0(\processor/wb_csr_data [25]),
        .I1(\csr_data_out[30]_i_8_n_0 ),
        .I2(\processor/csr_read_data [25]),
        .I3(\csr_data_out[30]_i_9_n_0 ),
        .I4(\processor/wb_exception_context[badaddr] [25]),
        .I5(\csr_data_out[4]_i_9_n_0 ),
        .O(\csr_data_out[25]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[26]_i_1 
       (.I0(\processor/ex_pc [26]),
        .I1(\processor/execute/csr_alu_instance/b [26]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[26]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[26]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[26]_i_2 
       (.I0(\processor/execute/rs1_forwarded [26]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FF07FF07FF07)) 
    \csr_data_out[26]_i_3 
       (.I0(\csr_data_out[30]_i_5_n_0 ),
        .I1(\processor/mem_csr_data [26]),
        .I2(\csr_data_out[26]_i_5_n_0 ),
        .I3(\csr_data_out[31]_i_6_n_0 ),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\processor/mem_exception_context[badaddr] [26]),
        .O(\csr_data_out[26]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[26]_i_4 
       (.I0(\processor/mem_rd_data [26]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [26]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [26]),
        .O(\processor/execute/rs1_forwarded [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFD800D8)) 
    \csr_data_out[26]_i_5 
       (.I0(\csr_data_out[30]_i_8_n_0 ),
        .I1(\processor/wb_csr_data [26]),
        .I2(\processor/csr_read_data [26]),
        .I3(\csr_data_out[30]_i_9_n_0 ),
        .I4(\processor/wb_exception_context[badaddr] [26]),
        .I5(\csr_data_out[4]_i_9_n_0 ),
        .O(\csr_data_out[26]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[27]_i_1 
       (.I0(\processor/ex_pc [27]),
        .I1(\processor/execute/csr_alu_instance/b [27]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[27]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[27]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[27]_i_2 
       (.I0(\processor/execute/rs1_forwarded [27]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FF07FF07FF07)) 
    \csr_data_out[27]_i_3 
       (.I0(\csr_data_out[30]_i_5_n_0 ),
        .I1(\processor/mem_csr_data [27]),
        .I2(\csr_data_out[27]_i_5_n_0 ),
        .I3(\csr_data_out[31]_i_6_n_0 ),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\processor/mem_exception_context[badaddr] [27]),
        .O(\csr_data_out[27]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[27]_i_4 
       (.I0(\processor/mem_rd_data [27]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [27]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [27]),
        .O(\processor/execute/rs1_forwarded [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFD800D8)) 
    \csr_data_out[27]_i_5 
       (.I0(\csr_data_out[30]_i_8_n_0 ),
        .I1(\processor/wb_csr_data [27]),
        .I2(\processor/csr_read_data [27]),
        .I3(\csr_data_out[30]_i_9_n_0 ),
        .I4(\processor/wb_exception_context[badaddr] [27]),
        .I5(\csr_data_out[4]_i_9_n_0 ),
        .O(\csr_data_out[27]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[28]_i_1 
       (.I0(\processor/ex_pc [28]),
        .I1(\processor/execute/csr_alu_instance/b [28]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[28]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[28]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[28]_i_2 
       (.I0(\processor/execute/rs1_forwarded [28]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FF07FF07FF07)) 
    \csr_data_out[28]_i_3 
       (.I0(\csr_data_out[30]_i_5_n_0 ),
        .I1(\processor/mem_csr_data [28]),
        .I2(\csr_data_out[28]_i_5_n_0 ),
        .I3(\csr_data_out[31]_i_6_n_0 ),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\processor/mem_exception_context[badaddr] [28]),
        .O(\csr_data_out[28]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[28]_i_4 
       (.I0(\processor/mem_rd_data [28]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [28]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [28]),
        .O(\processor/execute/rs1_forwarded [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFD800D8)) 
    \csr_data_out[28]_i_5 
       (.I0(\csr_data_out[30]_i_8_n_0 ),
        .I1(\processor/wb_csr_data [28]),
        .I2(\processor/csr_read_data [28]),
        .I3(\csr_data_out[30]_i_9_n_0 ),
        .I4(\processor/wb_exception_context[badaddr] [28]),
        .I5(\csr_data_out[4]_i_9_n_0 ),
        .O(\csr_data_out[28]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[29]_i_1 
       (.I0(\processor/ex_pc [29]),
        .I1(\processor/execute/csr_alu_instance/b [29]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[29]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[29]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[29]_i_2 
       (.I0(\processor/execute/rs1_forwarded [29]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FF07FF07FF07)) 
    \csr_data_out[29]_i_3 
       (.I0(\csr_data_out[30]_i_5_n_0 ),
        .I1(\processor/mem_csr_data [29]),
        .I2(\csr_data_out[29]_i_5_n_0 ),
        .I3(\csr_data_out[31]_i_6_n_0 ),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\processor/mem_exception_context[badaddr] [29]),
        .O(\csr_data_out[29]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[29]_i_4 
       (.I0(\processor/mem_rd_data [29]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [29]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [29]),
        .O(\processor/execute/rs1_forwarded [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    \csr_data_out[29]_i_5 
       (.I0(\processor/wb_csr_data [29]),
        .I1(\csr_data_out[30]_i_8_n_0 ),
        .I2(\processor/csr_read_data [29]),
        .I3(\csr_data_out[30]_i_9_n_0 ),
        .I4(\processor/wb_exception_context[badaddr] [29]),
        .I5(\csr_data_out[4]_i_9_n_0 ),
        .O(\csr_data_out[29]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[2]_i_1 
       (.I0(\processor/ex_pc [2]),
        .I1(\processor/execute/csr_alu_instance/b [2]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[2]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \csr_data_out[2]_i_2 
       (.I0(\processor/execute/rs1_addr [2]),
        .I1(\processor/execute/rs1_forwarded [2]),
        .I2(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000EEEEEEEF)) 
    \csr_data_out[2]_i_3 
       (.I0(\csr_data_out[2]_i_5_n_0 ),
        .I1(\csr_data_out[2]_i_6_n_0 ),
        .I2(\csr_data_out[2]_i_7_n_0 ),
        .I3(\csr_data_out[2]_i_8_n_0 ),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\csr_data_out[2]_i_9_n_0 ),
        .O(\csr_data_out[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[2]_i_4 
       (.I0(\processor/mem_rd_data [2]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [2]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [2]),
        .O(\processor/execute/rs1_forwarded [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000455500000000)) 
    \csr_data_out[2]_i_5 
       (.I0(\processor/wb_exception_context[cause] [2]),
        .I1(\csr_data_out[31]_i_18_n_0 ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/execute/csr_writeable ),
        .I4(\csr_data_out[31]_i_23_n_0 ),
        .I5(\processor/wb_exception ),
        .O(\csr_data_out[2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBAAAAAAAAAAAAA)) 
    \csr_data_out[2]_i_6 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\processor/mem_csr_data [2]),
        .I2(\processor/mem_csr_write [1]),
        .I3(\processor/mem_csr_write [0]),
        .I4(\processor/execute/csr_value_forwarded30_out ),
        .I5(\processor/execute/csr_writeable ),
        .O(\csr_data_out[2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[2]_i_7 
       (.I0(\processor/wb_exception_context[badaddr] [2]),
        .I1(\csr_data_out[31]_i_21_n_0 ),
        .O(\csr_data_out[2]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA888888808888888)) 
    \csr_data_out[2]_i_8 
       (.I0(\csr_data_out[31]_i_21_n_0 ),
        .I1(\processor/csr_read_data [2]),
        .I2(\processor/csr_unit/tohost_data1__0 ),
        .I3(\processor/execute/csr_value_forwarded3 ),
        .I4(\processor/execute/csr_writeable ),
        .I5(\processor/wb_csr_data [2]),
        .O(\csr_data_out[2]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \csr_data_out[2]_i_9 
       (.I0(\csr_data_out[31]_i_24_n_0 ),
        .I1(\processor/mem_exception_context[cause] [2]),
        .I2(\processor/mem_exception_context[badaddr] [2]),
        .I3(\csr_data_out[31]_i_25_n_0 ),
        .I4(\csr_data_out[4]_i_11_n_0 ),
        .O(\csr_data_out[2]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[30]_i_1 
       (.I0(\processor/ex_pc [30]),
        .I1(\processor/execute/csr_alu_instance/b [30]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[30]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[30]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFEFFFFFFFFFFFF)) 
    \csr_data_out[30]_i_10 
       (.I0(\processor/ex_csr_address[3]_repN ),
        .I1(\processor/ex_csr_address [5]),
        .I2(\csr_data_out[30]_i_11_n_0 ),
        .I3(\processor/ex_csr_address [4]),
        .I4(\processor/ex_csr_address [8]),
        .I5(\processor/ex_csr_address [9]),
        .O(\csr_data_out[30]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \csr_data_out[30]_i_11 
       (.I0(\processor/ex_csr_address [10]),
        .I1(\processor/ex_csr_address [11]),
        .I2(\processor/ex_csr_address [2]),
        .I3(\processor/ex_csr_address [7]),
        .O(\csr_data_out[30]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[30]_i_2 
       (.I0(\processor/execute/rs1_forwarded [30]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FF07FF07FF07)) 
    \csr_data_out[30]_i_3 
       (.I0(\csr_data_out[30]_i_5_n_0 ),
        .I1(\processor/mem_csr_data [30]),
        .I2(\csr_data_out[30]_i_6_n_0 ),
        .I3(\csr_data_out[31]_i_6_n_0 ),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\processor/mem_exception_context[badaddr] [30]),
        .O(\csr_data_out[30]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[30]_i_4 
       (.I0(\processor/mem_rd_data [30]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [30]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [30]),
        .O(\processor/execute/rs1_forwarded [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE000)) 
    \csr_data_out[30]_i_5 
       (.I0(\processor/mem_csr_write [1]),
        .I1(\processor/mem_csr_write [0]),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/execute/csr_writeable ),
        .O(\csr_data_out[30]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "csr_data_out[30]_i_5" *) 
  LUT4 #(
    .INIT(16'hE000)) 
    \csr_data_out[30]_i_5_replica 
       (.I0(\processor/mem_csr_write [1]),
        .I1(\processor/mem_csr_write [0]),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/execute/csr_writeable ),
        .O(\csr_data_out[30]_i_5_n_0_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFD800D8)) 
    \csr_data_out[30]_i_6 
       (.I0(\csr_data_out[30]_i_8_n_0 ),
        .I1(\processor/wb_csr_data [30]),
        .I2(\processor/csr_read_data [30]),
        .I3(\csr_data_out[30]_i_9_n_0 ),
        .I4(\processor/wb_exception_context[badaddr] [30]),
        .I5(\csr_data_out[4]_i_9_n_0 ),
        .O(\csr_data_out[30]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    \csr_data_out[30]_i_7 
       (.I0(\processor/mem_exception ),
        .I1(\processor/ex_csr_address [0]),
        .I2(\processor/ex_csr_address [1]),
        .I3(\processor/ex_csr_address[6]_repN ),
        .I4(\csr_data_out[31]_i_15_n_0 ),
        .I5(\csr_data_out[31]_i_14_n_0 ),
        .O(\csr_data_out[30]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8880)) 
    \csr_data_out[30]_i_8 
       (.I0(\processor/execute/csr_writeable ),
        .I1(\processor/execute/csr_value_forwarded3 ),
        .I2(\processor/wb_csr_write [1]),
        .I3(\processor/wb_csr_write [0]),
        .O(\csr_data_out[30]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00008000)) 
    \csr_data_out[30]_i_9 
       (.I0(\processor/wb_exception ),
        .I1(\processor/ex_csr_address [0]),
        .I2(\processor/ex_csr_address [1]),
        .I3(\processor/ex_csr_address[6]_repN ),
        .I4(\csr_data_out[30]_i_10_n_0 ),
        .O(\csr_data_out[30]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h4)) 
    \csr_data_out[31]_i_1 
       (.I0(reset),
        .I1(\processor/memory/p_1_in ),
        .O(\csr_data_out[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000A000CCCCACCC)) 
    \csr_data_out[31]_i_10 
       (.I0(\processor/mem_csr_data [31]),
        .I1(\csr_data_out[31]_i_16_n_0 ),
        .I2(\processor/execute/csr_writeable ),
        .I3(\processor/execute/csr_value_forwarded30_out ),
        .I4(\csr_data_out[31]_i_18_n_0 ),
        .I5(\csr_data_out[31]_i_19_n_0 ),
        .O(\csr_data_out[31]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4F44)) 
    \csr_data_out[31]_i_11 
       (.I0(\csr_data_out[31]_i_24_n_0 ),
        .I1(\processor/mem_exception_context[cause] [5]),
        .I2(\csr_data_out[31]_i_25_n_0 ),
        .I3(\processor/mem_exception_context[badaddr] [31]),
        .O(\csr_data_out[31]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000900900000000)) 
    \csr_data_out[31]_i_12 
       (.I0(\processor/mem_rd_address [3]),
        .I1(\processor/execute/rs1_addr [3]),
        .I2(\processor/execute/rs1_addr [4]),
        .I3(\processor/mem_rd_address [4]),
        .I4(registers_reg_r1_0_31_0_5_i_14_n_0),
        .I5(\dmem_data_out_p[31]_i_4_n_0 ),
        .O(\csr_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDFFDFFFFFFFFDFFD)) 
    \csr_data_out[31]_i_13 
       (.I0(\dmem_data_out_p[31]_i_6_n_0 ),
        .I1(\csr_data_out[31]_i_26_n_0 ),
        .I2(\processor/execute/rs1_addr [3]),
        .I3(\processor/wb_rd_address [3]),
        .I4(\processor/execute/rs1_addr [2]),
        .I5(\processor/wb_rd_address [2]),
        .O(\csr_data_out[31]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \csr_data_out[31]_i_14 
       (.I0(\processor/ex_csr_address [5]),
        .I1(\processor/ex_csr_address [2]),
        .I2(\processor/ex_csr_address [11]),
        .O(\csr_data_out[31]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFEFFFFFFFFFFFF)) 
    \csr_data_out[31]_i_15 
       (.I0(\processor/ex_csr_address[7]_repN ),
        .I1(\processor/ex_csr_address [10]),
        .I2(\processor/ex_csr_address [4]),
        .I3(\processor/ex_csr_address[3]_repN ),
        .I4(\processor/ex_csr_address [9]),
        .I5(\processor/ex_csr_address [8]),
        .O(\csr_data_out[31]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFF7FFFFFFFF)) 
    \csr_data_out[31]_i_16 
       (.I0(\processor/ex_csr_address [1]),
        .I1(\processor/ex_csr_address[6]_repN ),
        .I2(\csr_data_out[31]_i_15_n_0 ),
        .I3(\csr_data_out[31]_i_14_n_0 ),
        .I4(\processor/ex_csr_address [0]),
        .I5(\processor/wb_exception ),
        .O(\csr_data_out[31]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \csr_data_out[31]_i_18 
       (.I0(\processor/mem_csr_write [0]),
        .I1(\processor/mem_csr_write [1]),
        .O(\csr_data_out[31]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \csr_data_out[31]_i_19 
       (.I0(\processor/wb_exception ),
        .I1(\csr_data_out[11]_i_8_n_0 ),
        .I2(\processor/ex_csr_address [11]),
        .I3(\processor/ex_csr_address [2]),
        .I4(\processor/ex_csr_address [5]),
        .I5(\csr_data_out[31]_i_15_n_0 ),
        .O(\csr_data_out[31]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[31]_i_2 
       (.I0(\processor/ex_pc [31]),
        .I1(\processor/execute/csr_alu_instance/b [31]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[31]_i_4_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \csr_data_out[31]_i_20 
       (.I0(\processor/wb_exception_context[badaddr] [31]),
        .I1(\processor/wb_exception ),
        .I2(\csr_data_out[31]_i_14_n_0 ),
        .I3(\csr_data_out[31]_i_15_n_0 ),
        .I4(\csr_data_out[31]_i_31_n_0 ),
        .I5(\processor/ex_csr_address [0]),
        .O(\csr_data_out[31]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFF7FFFFFFFFF)) 
    \csr_data_out[31]_i_21 
       (.I0(\processor/ex_csr_address [0]),
        .I1(\processor/ex_csr_address [1]),
        .I2(\processor/ex_csr_address[6]_repN ),
        .I3(\csr_data_out[31]_i_15_n_0 ),
        .I4(\csr_data_out[31]_i_14_n_0 ),
        .I5(\processor/wb_exception ),
        .O(\csr_data_out[31]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \csr_data_out[31]_i_23 
       (.I0(\processor/ex_csr_address [0]),
        .I1(\processor/ex_csr_address [11]),
        .I2(\processor/ex_csr_address [2]),
        .I3(\processor/ex_csr_address [5]),
        .I4(\csr_data_out[31]_i_15_n_0 ),
        .I5(\csr_data_out[31]_i_31_n_0 ),
        .O(\csr_data_out[31]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFEFFFFFFFFFF)) 
    \csr_data_out[31]_i_24 
       (.I0(\csr_data_out[31]_i_31_n_0 ),
        .I1(\csr_data_out[31]_i_36_n_0 ),
        .I2(\csr_data_out[31]_i_37_n_0 ),
        .I3(\processor/ex_csr_address [8]),
        .I4(\processor/ex_csr_address [0]),
        .I5(\processor/mem_exception ),
        .O(\csr_data_out[31]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFDFFFFFFFFFFFF)) 
    \csr_data_out[31]_i_25 
       (.I0(\processor/ex_csr_address [0]),
        .I1(\csr_data_out[31]_i_31_n_0 ),
        .I2(\csr_data_out[31]_i_36_n_0 ),
        .I3(\csr_data_out[31]_i_37_n_0 ),
        .I4(\processor/ex_csr_address [8]),
        .I5(\processor/mem_exception ),
        .O(\csr_data_out[31]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    \csr_data_out[31]_i_26 
       (.I0(\processor/execute/rs1_addr [4]),
        .I1(\processor/wb_rd_address [4]),
        .I2(\processor/wb_rd_address [0]),
        .I3(\processor/execute/rs1_addr [0]),
        .I4(\processor/wb_rd_address [1]),
        .I5(\processor/execute/rs1_addr [1]),
        .O(\csr_data_out[31]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \csr_data_out[31]_i_27 
       (.I0(\processor/mem_csr_address [11]),
        .I1(\processor/ex_csr_address [11]),
        .I2(\processor/mem_csr_address [9]),
        .I3(\processor/ex_csr_address [9]),
        .I4(\processor/ex_csr_address [10]),
        .I5(\processor/mem_csr_address [10]),
        .O(\csr_data_out[31]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \csr_data_out[31]_i_28 
       (.I0(\processor/mem_csr_address [8]),
        .I1(\processor/ex_csr_address [8]),
        .I2(\processor/mem_csr_address [6]),
        .I3(\processor/ex_csr_address[6]_repN ),
        .I4(\processor/ex_csr_address[7]_repN ),
        .I5(\processor/mem_csr_address [7]),
        .O(\csr_data_out[31]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \csr_data_out[31]_i_29 
       (.I0(\processor/mem_csr_address [5]),
        .I1(\processor/ex_csr_address [5]),
        .I2(\processor/mem_csr_address[4]_repN ),
        .I3(\processor/ex_csr_address [4]),
        .I4(\processor/ex_csr_address[3]_repN ),
        .I5(\processor/mem_csr_address [3]),
        .O(\csr_data_out[31]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[31]_i_3 
       (.I0(\processor/execute/rs1_forwarded [31]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \csr_data_out[31]_i_30 
       (.I0(\processor/mem_csr_address [2]),
        .I1(\processor/ex_csr_address [2]),
        .I2(\processor/mem_csr_address [0]),
        .I3(\processor/ex_csr_address [0]),
        .I4(\processor/ex_csr_address [1]),
        .I5(\processor/mem_csr_address [1]),
        .O(\csr_data_out[31]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \csr_data_out[31]_i_31 
       (.I0(\processor/ex_csr_address[6]_repN ),
        .I1(\processor/ex_csr_address [1]),
        .O(\csr_data_out[31]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \csr_data_out[31]_i_32 
       (.I0(\processor/wb_csr_address [10]),
        .I1(\processor/ex_csr_address [10]),
        .I2(\processor/wb_csr_address [9]),
        .I3(\processor/ex_csr_address [9]),
        .I4(\processor/ex_csr_address [11]),
        .I5(\processor/wb_csr_address [11]),
        .O(\csr_data_out[31]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \csr_data_out[31]_i_33 
       (.I0(\processor/wb_csr_address [8]),
        .I1(\processor/ex_csr_address [8]),
        .I2(\processor/wb_csr_address [6]),
        .I3(\processor/ex_csr_address[6]_repN ),
        .I4(\processor/ex_csr_address[7]_repN ),
        .I5(\processor/wb_csr_address [7]),
        .O(\csr_data_out[31]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \csr_data_out[31]_i_34 
       (.I0(\processor/wb_csr_address [5]),
        .I1(\processor/ex_csr_address [5]),
        .I2(\processor/wb_csr_address [4]),
        .I3(\processor/ex_csr_address [4]),
        .I4(\processor/ex_csr_address[3]_repN ),
        .I5(\processor/wb_csr_address [3]),
        .O(\csr_data_out[31]_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \csr_data_out[31]_i_35 
       (.I0(\processor/wb_csr_address [2]),
        .I1(\processor/ex_csr_address [2]),
        .I2(\processor/wb_csr_address [0]),
        .I3(\processor/ex_csr_address [0]),
        .I4(\processor/ex_csr_address [1]),
        .I5(\processor/wb_csr_address [1]),
        .O(\csr_data_out[31]_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFD)) 
    \csr_data_out[31]_i_36 
       (.I0(\processor/ex_csr_address [9]),
        .I1(\processor/ex_csr_address [4]),
        .I2(\processor/ex_csr_address [5]),
        .I3(\processor/ex_csr_address[7]_repN ),
        .O(\csr_data_out[31]_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \csr_data_out[31]_i_37 
       (.I0(\processor/ex_csr_address [10]),
        .I1(\processor/ex_csr_address [11]),
        .I2(\processor/ex_csr_address [2]),
        .I3(\processor/ex_csr_address [3]),
        .O(\csr_data_out[31]_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000BABAFFBA)) 
    \csr_data_out[31]_i_4 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\csr_data_out[31]_i_7_n_0 ),
        .I2(\csr_data_out[31]_i_8_n_0 ),
        .I3(\csr_data_out[31]_i_9_n_0 ),
        .I4(\csr_data_out[31]_i_10_n_0 ),
        .I5(\csr_data_out[31]_i_11_n_0 ),
        .O(\csr_data_out[31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[31]_i_5 
       (.I0(\processor/mem_rd_data [31]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [31]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [31]),
        .O(\processor/execute/rs1_forwarded [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000008802)) 
    \csr_data_out[31]_i_6 
       (.I0(\processor/mem_exception ),
        .I1(\processor/ex_csr_address[6]_repN ),
        .I2(\processor/ex_csr_address [0]),
        .I3(\processor/ex_csr_address [1]),
        .I4(\csr_data_out[31]_i_14_n_0 ),
        .I5(\csr_data_out[31]_i_15_n_0 ),
        .O(\csr_data_out[31]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF55D5)) 
    \csr_data_out[31]_i_7 
       (.I0(\csr_data_out[31]_i_16_n_0 ),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\csr_data_out[31]_i_18_n_0 ),
        .I4(\csr_data_out[31]_i_19_n_0 ),
        .I5(\csr_data_out[31]_i_20_n_0 ),
        .O(\csr_data_out[31]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5555D5557FFFFFFF)) 
    \csr_data_out[31]_i_8 
       (.I0(\csr_data_out[31]_i_21_n_0 ),
        .I1(\processor/csr_unit/tohost_data1__0 ),
        .I2(\processor/execute/csr_value_forwarded3 ),
        .I3(\processor/execute/csr_writeable ),
        .I4(\processor/wb_csr_data [31]),
        .I5(\processor/csr_read_data [31]),
        .O(\csr_data_out[31]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF40FFFFFFFFFFFF)) 
    \csr_data_out[31]_i_9 
       (.I0(\csr_data_out[31]_i_18_n_0 ),
        .I1(\processor/execute/csr_value_forwarded30_out ),
        .I2(\processor/execute/csr_writeable ),
        .I3(\csr_data_out[31]_i_23_n_0 ),
        .I4(\processor/wb_exception ),
        .I5(\processor/wb_exception_context[cause] [5]),
        .O(\csr_data_out[31]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[3]_i_1 
       (.I0(\processor/ex_pc [3]),
        .I1(\processor/execute/csr_alu_instance/b [3]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[3]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    \csr_data_out[3]_i_10 
       (.I0(\csr_data_out[31]_i_31_n_0 ),
        .I1(\csr_data_out[3]_i_11_n_0 ),
        .I2(\csr_data_out[30]_i_11_n_0 ),
        .I3(\csr_data_out[3]_i_12_n_0 ),
        .I4(\processor/ex_csr_address [0]),
        .I5(\processor/wb_exception ),
        .O(\csr_data_out[3]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \csr_data_out[3]_i_11 
       (.I0(\processor/ex_csr_address [4]),
        .I1(\processor/ex_csr_address [8]),
        .I2(\processor/ex_csr_address [9]),
        .O(\csr_data_out[3]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \csr_data_out[3]_i_12 
       (.I0(\processor/ex_csr_address [5]),
        .I1(\processor/ex_csr_address [3]),
        .O(\csr_data_out[3]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \csr_data_out[3]_i_2 
       (.I0(\processor/execute/rs1_addr [3]),
        .I1(\processor/execute/rs1_forwarded [3]),
        .I2(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00FE)) 
    \csr_data_out[3]_i_3 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\csr_data_out[3]_i_5_n_0 ),
        .I2(\csr_data_out[3]_i_6_n_0 ),
        .I3(\csr_data_out[3]_i_7_n_0 ),
        .O(\csr_data_out[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[3]_i_4 
       (.I0(\processor/mem_rd_data [3]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [3]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [3]),
        .O(\processor/execute/rs1_forwarded [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000474700FF)) 
    \csr_data_out[3]_i_5 
       (.I0(\processor/wb_csr_data [3]),
        .I1(\csr_data_out[30]_i_8_n_0 ),
        .I2(\processor/csr_read_data [3]),
        .I3(\processor/wb_exception_context[badaddr] [3]),
        .I4(\csr_data_out[31]_i_21_n_0 ),
        .I5(\csr_data_out[4]_i_9_n_0 ),
        .O(\csr_data_out[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0070007000000070)) 
    \csr_data_out[3]_i_6 
       (.I0(\processor/mem_csr_data [3]),
        .I1(\csr_data_out[30]_i_5_n_0 ),
        .I2(\csr_data_out[4]_i_9_n_0 ),
        .I3(\csr_data_out[3]_i_8_n_0 ),
        .I4(\processor/wb_exception_context ),
        .I5(\csr_data_out[3]_i_9_n_0 ),
        .O(\csr_data_out[3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF44F444F444F4)) 
    \csr_data_out[3]_i_7 
       (.I0(\csr_data_out[31]_i_24_n_0 ),
        .I1(\processor/mem_exception_context[cause] [3]),
        .I2(\processor/mem_exception_context[badaddr] [3]),
        .I3(\csr_data_out[31]_i_25_n_0 ),
        .I4(\processor/mem_exception_context ),
        .I5(\csr_data_out[4]_i_11_n_0 ),
        .O(\csr_data_out[3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000001FFF0000)) 
    \csr_data_out[3]_i_8 
       (.I0(\processor/mem_csr_write [1]),
        .I1(\processor/mem_csr_write [0]),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/execute/csr_writeable ),
        .I4(\processor/wb_exception_context[cause] [3]),
        .I5(\csr_data_out[3]_i_10_n_0 ),
        .O(\csr_data_out[3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF08FF)) 
    \csr_data_out[3]_i_9 
       (.I0(\processor/execute/csr_writeable ),
        .I1(\processor/execute/csr_value_forwarded30_out ),
        .I2(\csr_data_out[31]_i_18_n_0 ),
        .I3(\processor/wb_exception ),
        .I4(\csr_data_out[11]_i_8_n_0 ),
        .I5(\csr_data_out[30]_i_10_n_0 ),
        .O(\csr_data_out[3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[4]_i_1 
       (.I0(\processor/ex_pc [4]),
        .I1(\processor/execute/csr_alu_instance/b [4]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[4]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \csr_data_out[4]_i_10 
       (.I0(\csr_data_out[31]_i_24_n_0 ),
        .I1(\processor/mem_exception_context[cause] [4]),
        .I2(\processor/mem_exception_context[badaddr] [4]),
        .I3(\csr_data_out[31]_i_25_n_0 ),
        .I4(\csr_data_out[4]_i_11_n_0 ),
        .O(\csr_data_out[4]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000020)) 
    \csr_data_out[4]_i_11 
       (.I0(\processor/mem_exception ),
        .I1(\csr_data_out[11]_i_8_n_0 ),
        .I2(\processor/ex_csr_address [8]),
        .I3(\csr_data_out[31]_i_37_n_0 ),
        .I4(\csr_data_out[31]_i_36_n_0 ),
        .O(\csr_data_out[4]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \csr_data_out[4]_i_2 
       (.I0(\processor/execute/rs1_addr [4]),
        .I1(\processor/execute/rs1_forwarded [4]),
        .I2(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000EEEEEEEF)) 
    \csr_data_out[4]_i_3 
       (.I0(\csr_data_out[4]_i_5_n_0 ),
        .I1(\csr_data_out[4]_i_6_n_0 ),
        .I2(\csr_data_out[4]_i_7_n_0 ),
        .I3(\csr_data_out[4]_i_8_n_0 ),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\csr_data_out[4]_i_10_n_0 ),
        .O(\csr_data_out[4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[4]_i_4 
       (.I0(\processor/mem_rd_data [4]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [4]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [4]),
        .O(\processor/execute/rs1_forwarded [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000455500000000)) 
    \csr_data_out[4]_i_5 
       (.I0(\processor/wb_exception_context[cause] [4]),
        .I1(\csr_data_out[31]_i_18_n_0 ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/execute/csr_writeable ),
        .I4(\csr_data_out[31]_i_23_n_0 ),
        .I5(\processor/wb_exception ),
        .O(\csr_data_out[4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBAAAAAAAAAAAAA)) 
    \csr_data_out[4]_i_6 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\processor/mem_csr_data [4]),
        .I2(\processor/mem_csr_write [1]),
        .I3(\processor/mem_csr_write [0]),
        .I4(\processor/execute/csr_value_forwarded30_out ),
        .I5(\processor/execute/csr_writeable ),
        .O(\csr_data_out[4]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[4]_i_7 
       (.I0(\processor/wb_exception_context[badaddr] [4]),
        .I1(\csr_data_out[31]_i_21_n_0 ),
        .O(\csr_data_out[4]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA888888808888888)) 
    \csr_data_out[4]_i_8 
       (.I0(\csr_data_out[31]_i_21_n_0 ),
        .I1(\processor/csr_read_data [4]),
        .I2(\processor/csr_unit/tohost_data1__0 ),
        .I3(\processor/execute/csr_value_forwarded3 ),
        .I4(\processor/execute/csr_writeable ),
        .I5(\processor/wb_csr_data [4]),
        .O(\csr_data_out[4]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBAAABAAAFFFFBAAA)) 
    \csr_data_out[4]_i_9 
       (.I0(\csr_data_out[31]_i_19_n_0 ),
        .I1(\csr_data_out[31]_i_18_n_0 ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/execute/csr_writeable ),
        .I4(\processor/wb_exception ),
        .I5(\csr_data_out[31]_i_23_n_0 ),
        .O(\csr_data_out[4]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[5]_i_1 
       (.I0(\processor/ex_pc [5]),
        .I1(\processor/execute/csr_alu_instance/b [5]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[5]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[5]_i_2 
       (.I0(\processor/execute/rs1_forwarded [5]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000F2F2F2)) 
    \csr_data_out[5]_i_3 
       (.I0(\csr_data_out[5]_i_5_n_0 ),
        .I1(\csr_data_out[5]_i_6_n_0 ),
        .I2(\csr_data_out[31]_i_6_n_0 ),
        .I3(\processor/mem_exception_context[badaddr] [5]),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\csr_data_out[11]_i_7_n_0 ),
        .O(\csr_data_out[5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[5]_i_4 
       (.I0(\processor/mem_rd_data [5]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [5]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [5]),
        .O(\processor/execute/rs1_forwarded [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAABABFFFFFBABF)) 
    \csr_data_out[5]_i_5 
       (.I0(\csr_data_out[4]_i_9_n_0 ),
        .I1(\processor/wb_csr_data [5]),
        .I2(\csr_data_out[30]_i_8_n_0 ),
        .I3(\processor/csr_read_data [5]),
        .I4(\csr_data_out[30]_i_9_n_0 ),
        .I5(\processor/wb_exception_context[badaddr] [5]),
        .O(\csr_data_out[5]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFFFFFFA8000000)) 
    \csr_data_out[5]_i_6 
       (.I0(\processor/mem_csr_data [5]),
        .I1(\processor/mem_csr_write [1]),
        .I2(\processor/mem_csr_write [0]),
        .I3(\processor/execute/csr_value_forwarded30_out ),
        .I4(\processor/execute/csr_writeable ),
        .I5(\csr_data_out[31]_i_19_n_0 ),
        .O(\csr_data_out[5]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[6]_i_1 
       (.I0(\processor/ex_pc [6]),
        .I1(\processor/execute/csr_alu_instance/b [6]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[6]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[6]_i_2 
       (.I0(\processor/execute/rs1_forwarded [6]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FF07FF07FF07)) 
    \csr_data_out[6]_i_3 
       (.I0(\csr_data_out[30]_i_5_n_0_repN ),
        .I1(\processor/mem_csr_data [6]),
        .I2(\csr_data_out[6]_i_5_n_0 ),
        .I3(\csr_data_out[31]_i_6_n_0 ),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\processor/mem_exception_context[badaddr] [6]),
        .O(\csr_data_out[6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[6]_i_4 
       (.I0(\processor/mem_rd_data [6]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [6]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [6]),
        .O(\processor/execute/rs1_forwarded [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    \csr_data_out[6]_i_5 
       (.I0(\processor/wb_csr_data [6]),
        .I1(\csr_data_out[30]_i_8_n_0 ),
        .I2(\processor/csr_read_data [6]),
        .I3(\csr_data_out[30]_i_9_n_0 ),
        .I4(\processor/wb_exception_context[badaddr] [6]),
        .I5(\csr_data_out[4]_i_9_n_0 ),
        .O(\csr_data_out[6]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[7]_i_1 
       (.I0(\processor/ex_pc [7]),
        .I1(\processor/execute/csr_alu_instance/b [7]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[7]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[7]_i_2 
       (.I0(\processor/execute/rs1_forwarded [7]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000F2F2F2)) 
    \csr_data_out[7]_i_3 
       (.I0(\csr_data_out[7]_i_5_n_0 ),
        .I1(\csr_data_out[7]_i_6_n_0 ),
        .I2(\csr_data_out[31]_i_6_n_0 ),
        .I3(\processor/mem_exception_context[badaddr] [7]),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\csr_data_out[11]_i_7_n_0 ),
        .O(\csr_data_out[7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[7]_i_4 
       (.I0(\processor/mem_rd_data[7]_repN_1 ),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [7]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [7]),
        .O(\processor/execute/rs1_forwarded [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "csr_data_out[7]_i_4" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[7]_i_4_replica 
       (.I0(\processor/mem_rd_data[7]_repN ),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [7]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [7]),
        .O(\processor/execute/rs1_forwarded[7]_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAABABFFFFFBABF)) 
    \csr_data_out[7]_i_5 
       (.I0(\csr_data_out[4]_i_9_n_0 ),
        .I1(\processor/wb_csr_data [7]),
        .I2(\csr_data_out[30]_i_8_n_0 ),
        .I3(\processor/csr_read_data [7]),
        .I4(\csr_data_out[30]_i_9_n_0 ),
        .I5(\processor/wb_exception_context[badaddr] [7]),
        .O(\csr_data_out[7]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFFFFFFA8000000)) 
    \csr_data_out[7]_i_6 
       (.I0(\processor/mem_csr_data [7]),
        .I1(\processor/mem_csr_write [1]),
        .I2(\processor/mem_csr_write [0]),
        .I3(\processor/execute/csr_value_forwarded30_out ),
        .I4(\processor/execute/csr_writeable ),
        .I5(\csr_data_out[31]_i_19_n_0 ),
        .O(\csr_data_out[7]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[8]_i_1 
       (.I0(\processor/ex_pc [8]),
        .I1(\processor/execute/csr_alu_instance/b [8]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[8]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[8]_i_2 
       (.I0(\processor/execute/rs1_forwarded [8]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000F2F2F2)) 
    \csr_data_out[8]_i_3 
       (.I0(\csr_data_out[8]_i_5_n_0 ),
        .I1(\csr_data_out[8]_i_6_n_0 ),
        .I2(\csr_data_out[31]_i_6_n_0 ),
        .I3(\processor/mem_exception_context[badaddr] [8]),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\csr_data_out[11]_i_7_n_0 ),
        .O(\csr_data_out[8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[8]_i_4 
       (.I0(\processor/mem_rd_data [8]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [8]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [8]),
        .O(\processor/execute/rs1_forwarded [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAABABFFFFFBABF)) 
    \csr_data_out[8]_i_5 
       (.I0(\csr_data_out[4]_i_9_n_0 ),
        .I1(\processor/wb_csr_data [8]),
        .I2(\csr_data_out[30]_i_8_n_0 ),
        .I3(\processor/csr_read_data [8]),
        .I4(\csr_data_out[30]_i_9_n_0 ),
        .I5(\processor/wb_exception_context[badaddr] [8]),
        .O(\csr_data_out[8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFFFFFFA8000000)) 
    \csr_data_out[8]_i_6 
       (.I0(\processor/mem_csr_data [8]),
        .I1(\processor/mem_csr_write [1]),
        .I2(\processor/mem_csr_write [0]),
        .I3(\processor/execute/csr_value_forwarded30_out ),
        .I4(\processor/execute/csr_writeable ),
        .I5(\csr_data_out[31]_i_19_n_0 ),
        .O(\csr_data_out[8]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAACCCF003F)) 
    \csr_data_out[9]_i_1 
       (.I0(\processor/ex_pc [9]),
        .I1(\processor/execute/csr_alu_instance/b [9]),
        .I2(\processor/ex_csr_write [1]),
        .I3(\csr_data_out[9]_i_3_n_0 ),
        .I4(\processor/ex_csr_write [0]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\csr_data_out[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \csr_data_out[9]_i_2 
       (.I0(\processor/execute/rs1_forwarded [9]),
        .I1(\processor/execute/funct3 [2]),
        .O(\processor/execute/csr_alu_instance/b [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FF07FF07FF07)) 
    \csr_data_out[9]_i_3 
       (.I0(\csr_data_out[30]_i_5_n_0 ),
        .I1(\processor/mem_csr_data [9]),
        .I2(\csr_data_out[9]_i_5_n_0 ),
        .I3(\csr_data_out[31]_i_6_n_0 ),
        .I4(\csr_data_out[30]_i_7_n_0 ),
        .I5(\processor/mem_exception_context[badaddr] [9]),
        .O(\csr_data_out[9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \csr_data_out[9]_i_4 
       (.I0(\processor/mem_rd_data [9]),
        .I1(\csr_data_out[31]_i_12_n_0 ),
        .I2(\processor/rs1_data [9]),
        .I3(\csr_data_out[31]_i_13_n_0 ),
        .I4(\processor/wb_rd_data [9]),
        .O(\processor/execute/rs1_forwarded [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFD800D8)) 
    \csr_data_out[9]_i_5 
       (.I0(\csr_data_out[30]_i_8_n_0 ),
        .I1(\processor/wb_csr_data [9]),
        .I2(\processor/csr_read_data [9]),
        .I3(\csr_data_out[30]_i_9_n_0 ),
        .I4(\processor/wb_exception_context[badaddr] [9]),
        .I5(\csr_data_out[4]_i_9_n_0 ),
        .O(\csr_data_out[9]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \csr_data_out_reg[31]_i_17 
       (.CI(\<const0>__0__0 ),
        .CO({\processor/execute/csr_value_forwarded30_out ,\csr_data_out_reg[31]_i_17_n_1 ,\csr_data_out_reg[31]_i_17_n_2 ,\csr_data_out_reg[31]_i_17_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\csr_data_out[31]_i_27_n_0 ,\csr_data_out[31]_i_28_n_0 ,\csr_data_out[31]_i_29_n_0 ,\csr_data_out[31]_i_30_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \csr_data_out_reg[31]_i_22 
       (.CI(\<const0>__0__0 ),
        .CO({\processor/execute/csr_value_forwarded3 ,\csr_data_out_reg[31]_i_22_n_1 ,\csr_data_out_reg[31]_i_22_n_2 ,\csr_data_out_reg[31]_i_22_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\csr_data_out[31]_i_32_n_0 ,\csr_data_out[31]_i_33_n_0 ,\csr_data_out[31]_i_34_n_0 ,\csr_data_out[31]_i_35_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAABAAAAAAAA)) 
    \csr_read_address_p[0]_i_1 
       (.I0(\processor/id_immediate [0]),
        .I1(\csr_read_address_p[0]_i_2_n_0 ),
        .I2(\csr_read_address_p[0]_i_3_n_0 ),
        .I3(\csr_read_address_p[0]_i_4_n_0 ),
        .I4(\csr_read_address_p[0]_i_5_n_0 ),
        .I5(\processor/id_immediate [8]),
        .O(\processor/decode/csr_addr__40 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFEF0F0)) 
    \csr_read_address_p[0]_i_2 
       (.I0(data0[26]),
        .I1(data0[27]),
        .I2(\processor/id_immediate [1]),
        .I3(data0[29]),
        .I4(\csr_addr[10]_i_2_n_0 ),
        .O(\csr_read_address_p[0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \csr_read_address_p[0]_i_3 
       (.I0(\processor/id_immediate [3]),
        .I1(\processor/id_immediate [2]),
        .O(\csr_read_address_p[0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF8)) 
    \csr_read_address_p[0]_i_4 
       (.I0(\csr_addr[10]_i_2_n_0 ),
        .I1(data0[25]),
        .I2(\processor/id_immediate [4]),
        .O(\csr_read_address_p[0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF8)) 
    \csr_read_address_p[0]_i_5 
       (.I0(\csr_addr[10]_i_2_n_0 ),
        .I1(data0[30]),
        .I2(\processor/id_immediate [11]),
        .O(\csr_read_address_p[0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h200020000000A02A)) 
    \csr_read_address_p[0]_i_6 
       (.I0(data0[28]),
        .I1(\processor/decode/instruction_reg_n_0_[4] ),
        .I2(\processor/decode/instruction_reg_n_0_[5] ),
        .I3(\processor/decode/instruction_reg_n_0_[6] ),
        .I4(\processor/decode/instruction_reg_n_0_[3] ),
        .I5(\processor/decode/instruction_reg_n_0_ ),
        .O(\processor/id_immediate [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h200020000000A02A)) 
    \csr_read_address_p[10]_i_1 
       (.I0(data0[30]),
        .I1(\processor/decode/instruction_reg_n_0_[4] ),
        .I2(\processor/decode/instruction_reg_n_0_[5] ),
        .I3(\processor/decode/instruction_reg_n_0_[6] ),
        .I4(\processor/decode/instruction_reg_n_0_[3] ),
        .I5(\processor/decode/instruction_reg_n_0_ ),
        .O(\processor/id_immediate [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h4)) 
    \csr_read_address_p[11]_i_1 
       (.I0(\csr_addr[11]_i_2_n_0 ),
        .I1(\processor/execute/exception_taken0 ),
        .O(\csr_read_address_p[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h200020000000A02A)) 
    \csr_read_address_p[5]_i_1 
       (.I0(data0[25]),
        .I1(\processor/decode/instruction_reg_n_0_[4] ),
        .I2(\processor/decode/instruction_reg_n_0_[5] ),
        .I3(\processor/decode/instruction_reg_n_0_[6] ),
        .I4(\processor/decode/instruction_reg_n_0_[3] ),
        .I5(\processor/decode/instruction_reg_n_0_ ),
        .O(\processor/id_immediate [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF8)) 
    \csr_read_address_p[6]_i_1 
       (.I0(\csr_addr[10]_i_2_n_0 ),
        .I1(data0[26]),
        .I2(\csr_addr[9]_i_2_n_0 ),
        .O(\processor/decode/csr_addr__40 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h200020000000A02A)) 
    \csr_read_address_p[7]_i_1 
       (.I0(data0[27]),
        .I1(\processor/decode/instruction_reg_n_0_[4] ),
        .I2(\processor/decode/instruction_reg_n_0_[5] ),
        .I3(\processor/decode/instruction_reg_n_0_[6] ),
        .I4(\processor/decode/instruction_reg_n_0_[3] ),
        .I5(\processor/decode/instruction_reg_n_0_ ),
        .O(\processor/id_immediate [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF8)) 
    \csr_read_address_p[8]_i_1 
       (.I0(\csr_addr[10]_i_2_n_0 ),
        .I1(data0[28]),
        .I2(\csr_addr[9]_i_2_n_0 ),
        .O(\processor/decode/csr_addr__40 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF8)) 
    \csr_read_address_p[9]_i_1 
       (.I0(\csr_addr[10]_i_2_n_0 ),
        .I1(data0[29]),
        .I2(\csr_addr[9]_i_2_n_0 ),
        .O(\processor/decode/csr_addr__40 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000101000)) 
    \csr_write[0]_i_1 
       (.I0(\processor/decode/instruction_reg_n_0_ ),
        .I1(\processor/decode/instruction_reg_n_0_[3] ),
        .I2(\processor/decode/instruction_reg_n_0_[6] ),
        .I3(\processor/id_funct3 [1]),
        .I4(\processor/id_funct3 [0]),
        .I5(csr_write),
        .O(\processor/id_csr_write [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \csr_write[0]_i_2 
       (.I0(\processor/decode/instruction_reg_n_0_[5] ),
        .I1(\processor/decode/instruction_reg_n_0_[4] ),
        .O(csr_write));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \csr_write[1]_i_1 
       (.I0(\processor/decode/instruction_reg_n_0_ ),
        .I1(\processor/decode/instruction_reg_n_0_[3] ),
        .I2(\processor/decode/instruction_reg_n_0_[6] ),
        .I3(\processor/id_funct3 [0]),
        .I4(\processor/decode/instruction_reg_n_0_[5] ),
        .I5(\processor/decode/instruction_reg_n_0_[4] ),
        .O(\processor/id_csr_write [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \csr_write_out[1]_i_1 
       (.I0(reset),
        .O(\icache/p_3_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFAFAFFCF)) 
    \csr_write_out[1]_i_2 
       (.I0(dmem_read_ack),
        .I1(dmem_write_ack),
        .I2(\processor/mem_mem_op [2]),
        .I3(\processor/mem_mem_op [0]),
        .I4(\processor/mem_mem_op [1]),
        .O(\processor/memory/p_1_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h10000000)) 
    \csr_write_out[1]_i_3 
       (.I0(\dmem_if/state_reg_n_0_ ),
        .I1(\arbiter/state [0]),
        .I2(wb_ack_in),
        .I3(\arbiter/state [1]),
        .I4(\dmem_if/state_reg_n_0_[1] ),
        .O(dmem_write_ack));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    csr_writeable_i_1
       (.I0(\csr_addr[11]_i_1_n_0 ),
        .I1(\csr_addr[10]_i_1_n_0 ),
        .O(\processor/csr_read_writeable ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \current_count[0]_i_5 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_ ),
        .O(\current_count[0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \current_count[0]_i_5__0 
       (.I0(\processor/csr_unit/cycle_counter/current_count_reg_n_0_ ),
        .O(current_count));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \current_count[0]_i_5__1 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_ ),
        .O(\current_count[0]_i_5__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[0]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO({\current_count_reg[0]_i_1_n_0 ,\current_count_reg[0]_i_1_n_1 ,\current_count_reg[0]_i_1_n_2 ,\current_count_reg[0]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .O({\current_count_reg[0]_i_1_n_4 ,\current_count_reg[0]_i_1_n_5 ,\current_count_reg[0]_i_1_n_6 ,\current_count_reg[0]_i_1_n_7 }),
        .S({\processor/csr_unit/timer_counter/current_count_reg_n_0_[3] ,\processor/csr_unit/timer_counter/current_count_reg_n_0_[2] ,\processor/csr_unit/timer_counter/current_count_reg_n_0_[1] ,\current_count[0]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[0]_i_1__0 
       (.CI(\<const0>__0__0 ),
        .CO(current_count_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .O({\current_count_reg[0]_i_1__0_n_4 ,\current_count_reg[0]_i_1__0_n_5 ,\current_count_reg[0]_i_1__0_n_6 ,\current_count_reg[0]_i_1__0_n_7 }),
        .S({\processor/csr_unit/cycle_counter/current_count_reg_n_0_[3] ,\processor/csr_unit/cycle_counter/current_count_reg_n_0_[2] ,\processor/csr_unit/cycle_counter/current_count_reg_n_0_[1] ,current_count}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[0]_i_1__1 
       (.CI(\<const0>__0__0 ),
        .CO({\current_count_reg[0]_i_1__1_n_0 ,\current_count_reg[0]_i_1__1_n_1 ,\current_count_reg[0]_i_1__1_n_2 ,\current_count_reg[0]_i_1__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .O({\current_count_reg[0]_i_1__1_n_4 ,\current_count_reg[0]_i_1__1_n_5 ,\current_count_reg[0]_i_1__1_n_6 ,\current_count_reg[0]_i_1__1_n_7 }),
        .S({\processor/csr_unit/instret_counter/current_count_reg_n_0_[3] ,\processor/csr_unit/instret_counter/current_count_reg_n_0_[2] ,\processor/csr_unit/instret_counter/current_count_reg_n_0_[1] ,\current_count[0]_i_5__1_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[12]_i_1 
       (.CI(\current_count_reg[8]_i_1_n_0 ),
        .CO({\current_count_reg[12]_i_1_n_0 ,\current_count_reg[12]_i_1_n_1 ,\current_count_reg[12]_i_1_n_2 ,\current_count_reg[12]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[12]_i_1_n_4 ,\current_count_reg[12]_i_1_n_5 ,\current_count_reg[12]_i_1_n_6 ,\current_count_reg[12]_i_1_n_7 }),
        .S({\processor/csr_unit/timer_counter/current_count_reg_n_0_[15] ,\processor/csr_unit/timer_counter/current_count_reg_n_0_[14] ,\processor/csr_unit/timer_counter/current_count_reg_n_0_[13] ,\processor/csr_unit/timer_counter/current_count_reg_n_0_[12] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[12]_i_1__0 
       (.CI(\current_count_reg[8]_i_1__0_n_0 ),
        .CO({\current_count_reg[12]_i_1__0_n_0 ,\current_count_reg[12]_i_1__0_n_1 ,\current_count_reg[12]_i_1__0_n_2 ,\current_count_reg[12]_i_1__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[12]_i_1__0_n_4 ,\current_count_reg[12]_i_1__0_n_5 ,\current_count_reg[12]_i_1__0_n_6 ,\current_count_reg[12]_i_1__0_n_7 }),
        .S({\processor/csr_unit/cycle_counter/current_count_reg_n_0_[15] ,\processor/csr_unit/cycle_counter/current_count_reg_n_0_[14] ,\processor/csr_unit/cycle_counter/current_count_reg_n_0_[13] ,\processor/csr_unit/cycle_counter/current_count_reg_n_0_[12] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[12]_i_1__1 
       (.CI(\current_count_reg[8]_i_1__1_n_0 ),
        .CO({\current_count_reg[12]_i_1__1_n_0 ,\current_count_reg[12]_i_1__1_n_1 ,\current_count_reg[12]_i_1__1_n_2 ,\current_count_reg[12]_i_1__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[12]_i_1__1_n_4 ,\current_count_reg[12]_i_1__1_n_5 ,\current_count_reg[12]_i_1__1_n_6 ,\current_count_reg[12]_i_1__1_n_7 }),
        .S({\processor/csr_unit/instret_counter/current_count_reg_n_0_[15] ,\processor/csr_unit/instret_counter/current_count_reg_n_0_[14] ,\processor/csr_unit/instret_counter/current_count_reg_n_0_[13] ,\processor/csr_unit/instret_counter/current_count_reg_n_0_[12] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[16]_i_1 
       (.CI(\current_count_reg[12]_i_1_n_0 ),
        .CO({\current_count_reg[16]_i_1_n_0 ,\current_count_reg[16]_i_1_n_1 ,\current_count_reg[16]_i_1_n_2 ,\current_count_reg[16]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[16]_i_1_n_4 ,\current_count_reg[16]_i_1_n_5 ,\current_count_reg[16]_i_1_n_6 ,\current_count_reg[16]_i_1_n_7 }),
        .S({\processor/csr_unit/timer_counter/current_count_reg_n_0_[19] ,\processor/csr_unit/timer_counter/current_count_reg_n_0_[18] ,\processor/csr_unit/timer_counter/current_count_reg_n_0_[17] ,\processor/csr_unit/timer_counter/current_count_reg_n_0_[16] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[16]_i_1__0 
       (.CI(\current_count_reg[12]_i_1__0_n_0 ),
        .CO({\current_count_reg[16]_i_1__0_n_0 ,\current_count_reg[16]_i_1__0_n_1 ,\current_count_reg[16]_i_1__0_n_2 ,\current_count_reg[16]_i_1__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[16]_i_1__0_n_4 ,\current_count_reg[16]_i_1__0_n_5 ,\current_count_reg[16]_i_1__0_n_6 ,\current_count_reg[16]_i_1__0_n_7 }),
        .S({\processor/csr_unit/cycle_counter/current_count_reg_n_0_[19] ,\processor/csr_unit/cycle_counter/current_count_reg_n_0_[18] ,\processor/csr_unit/cycle_counter/current_count_reg_n_0_[17] ,\processor/csr_unit/cycle_counter/current_count_reg_n_0_[16] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[16]_i_1__1 
       (.CI(\current_count_reg[12]_i_1__1_n_0 ),
        .CO({\current_count_reg[16]_i_1__1_n_0 ,\current_count_reg[16]_i_1__1_n_1 ,\current_count_reg[16]_i_1__1_n_2 ,\current_count_reg[16]_i_1__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[16]_i_1__1_n_4 ,\current_count_reg[16]_i_1__1_n_5 ,\current_count_reg[16]_i_1__1_n_6 ,\current_count_reg[16]_i_1__1_n_7 }),
        .S({\processor/csr_unit/instret_counter/current_count_reg_n_0_[19] ,\processor/csr_unit/instret_counter/current_count_reg_n_0_[18] ,\processor/csr_unit/instret_counter/current_count_reg_n_0_[17] ,\processor/csr_unit/instret_counter/current_count_reg_n_0_[16] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[20]_i_1 
       (.CI(\current_count_reg[16]_i_1_n_0 ),
        .CO({\current_count_reg[20]_i_1_n_0 ,\current_count_reg[20]_i_1_n_1 ,\current_count_reg[20]_i_1_n_2 ,\current_count_reg[20]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[20]_i_1_n_4 ,\current_count_reg[20]_i_1_n_5 ,\current_count_reg[20]_i_1_n_6 ,\current_count_reg[20]_i_1_n_7 }),
        .S({\processor/csr_unit/timer_counter/current_count_reg_n_0_[23] ,\processor/csr_unit/timer_counter/current_count_reg_n_0_[22] ,\processor/csr_unit/timer_counter/current_count_reg_n_0_[21] ,\processor/csr_unit/timer_counter/current_count_reg_n_0_[20] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[20]_i_1__0 
       (.CI(\current_count_reg[16]_i_1__0_n_0 ),
        .CO({\current_count_reg[20]_i_1__0_n_0 ,\current_count_reg[20]_i_1__0_n_1 ,\current_count_reg[20]_i_1__0_n_2 ,\current_count_reg[20]_i_1__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[20]_i_1__0_n_4 ,\current_count_reg[20]_i_1__0_n_5 ,\current_count_reg[20]_i_1__0_n_6 ,\current_count_reg[20]_i_1__0_n_7 }),
        .S({\processor/csr_unit/cycle_counter/current_count_reg_n_0_[23] ,\processor/csr_unit/cycle_counter/current_count_reg_n_0_[22] ,\processor/csr_unit/cycle_counter/current_count_reg_n_0_[21] ,\processor/csr_unit/cycle_counter/current_count_reg_n_0_[20] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[20]_i_1__1 
       (.CI(\current_count_reg[16]_i_1__1_n_0 ),
        .CO({\current_count_reg[20]_i_1__1_n_0 ,\current_count_reg[20]_i_1__1_n_1 ,\current_count_reg[20]_i_1__1_n_2 ,\current_count_reg[20]_i_1__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[20]_i_1__1_n_4 ,\current_count_reg[20]_i_1__1_n_5 ,\current_count_reg[20]_i_1__1_n_6 ,\current_count_reg[20]_i_1__1_n_7 }),
        .S({\processor/csr_unit/instret_counter/current_count_reg_n_0_[23] ,\processor/csr_unit/instret_counter/current_count_reg_n_0_[22] ,\processor/csr_unit/instret_counter/current_count_reg_n_0_[21] ,\processor/csr_unit/instret_counter/current_count_reg_n_0_[20] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[24]_i_1 
       (.CI(\current_count_reg[20]_i_1_n_0 ),
        .CO({\current_count_reg[24]_i_1_n_0 ,\current_count_reg[24]_i_1_n_1 ,\current_count_reg[24]_i_1_n_2 ,\current_count_reg[24]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[24]_i_1_n_4 ,\current_count_reg[24]_i_1_n_5 ,\current_count_reg[24]_i_1_n_6 ,\current_count_reg[24]_i_1_n_7 }),
        .S({\processor/csr_unit/timer_counter/current_count_reg_n_0_[27] ,\processor/csr_unit/timer_counter/current_count_reg_n_0_[26] ,\processor/csr_unit/timer_counter/current_count_reg_n_0_[25] ,\processor/csr_unit/timer_counter/current_count_reg_n_0_[24] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[24]_i_1__0 
       (.CI(\current_count_reg[20]_i_1__0_n_0 ),
        .CO({\current_count_reg[24]_i_1__0_n_0 ,\current_count_reg[24]_i_1__0_n_1 ,\current_count_reg[24]_i_1__0_n_2 ,\current_count_reg[24]_i_1__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[24]_i_1__0_n_4 ,\current_count_reg[24]_i_1__0_n_5 ,\current_count_reg[24]_i_1__0_n_6 ,\current_count_reg[24]_i_1__0_n_7 }),
        .S({\processor/csr_unit/cycle_counter/current_count_reg_n_0_[27] ,\processor/csr_unit/cycle_counter/current_count_reg_n_0_[26] ,\processor/csr_unit/cycle_counter/current_count_reg_n_0_[25] ,\processor/csr_unit/cycle_counter/current_count_reg_n_0_[24] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[24]_i_1__1 
       (.CI(\current_count_reg[20]_i_1__1_n_0 ),
        .CO({\current_count_reg[24]_i_1__1_n_0 ,\current_count_reg[24]_i_1__1_n_1 ,\current_count_reg[24]_i_1__1_n_2 ,\current_count_reg[24]_i_1__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[24]_i_1__1_n_4 ,\current_count_reg[24]_i_1__1_n_5 ,\current_count_reg[24]_i_1__1_n_6 ,\current_count_reg[24]_i_1__1_n_7 }),
        .S({\processor/csr_unit/instret_counter/current_count_reg_n_0_[27] ,\processor/csr_unit/instret_counter/current_count_reg_n_0_[26] ,\processor/csr_unit/instret_counter/current_count_reg_n_0_[25] ,\processor/csr_unit/instret_counter/current_count_reg_n_0_[24] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[28]_i_1 
       (.CI(\current_count_reg[24]_i_1_n_0 ),
        .CO({\current_count_reg[28]_i_1_n_0 ,\current_count_reg[28]_i_1_n_1 ,\current_count_reg[28]_i_1_n_2 ,\current_count_reg[28]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[28]_i_1_n_4 ,\current_count_reg[28]_i_1_n_5 ,\current_count_reg[28]_i_1_n_6 ,\current_count_reg[28]_i_1_n_7 }),
        .S({\processor/csr_unit/timer_counter/current_count_reg_n_0_[31] ,\processor/csr_unit/timer_counter/current_count_reg_n_0_[30] ,\processor/csr_unit/timer_counter/current_count_reg_n_0_[29] ,\processor/csr_unit/timer_counter/current_count_reg_n_0_[28] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[28]_i_1__0 
       (.CI(\current_count_reg[24]_i_1__0_n_0 ),
        .CO({\current_count_reg[28]_i_1__0_n_0 ,\current_count_reg[28]_i_1__0_n_1 ,\current_count_reg[28]_i_1__0_n_2 ,\current_count_reg[28]_i_1__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[28]_i_1__0_n_4 ,\current_count_reg[28]_i_1__0_n_5 ,\current_count_reg[28]_i_1__0_n_6 ,\current_count_reg[28]_i_1__0_n_7 }),
        .S({\processor/csr_unit/cycle_counter/current_count_reg_n_0_[31] ,\processor/csr_unit/cycle_counter/current_count_reg_n_0_[30] ,\processor/csr_unit/cycle_counter/current_count_reg_n_0_[29] ,\processor/csr_unit/cycle_counter/current_count_reg_n_0_[28] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[28]_i_1__1 
       (.CI(\current_count_reg[24]_i_1__1_n_0 ),
        .CO({\current_count_reg[28]_i_1__1_n_0 ,\current_count_reg[28]_i_1__1_n_1 ,\current_count_reg[28]_i_1__1_n_2 ,\current_count_reg[28]_i_1__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[28]_i_1__1_n_4 ,\current_count_reg[28]_i_1__1_n_5 ,\current_count_reg[28]_i_1__1_n_6 ,\current_count_reg[28]_i_1__1_n_7 }),
        .S({\processor/csr_unit/instret_counter/current_count_reg_n_0_[31] ,\processor/csr_unit/instret_counter/current_count_reg_n_0_[30] ,\processor/csr_unit/instret_counter/current_count_reg_n_0_[29] ,\processor/csr_unit/instret_counter/current_count_reg_n_0_[28] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[32]_i_1 
       (.CI(\current_count_reg[28]_i_1_n_0 ),
        .CO({\current_count_reg[32]_i_1_n_0 ,\current_count_reg[32]_i_1_n_1 ,\current_count_reg[32]_i_1_n_2 ,\current_count_reg[32]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[32]_i_1_n_4 ,\current_count_reg[32]_i_1_n_5 ,\current_count_reg[32]_i_1_n_6 ,\current_count_reg[32]_i_1_n_7 }),
        .S(data12[3:0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[32]_i_1__0 
       (.CI(\current_count_reg[28]_i_1__0_n_0 ),
        .CO({\current_count_reg[32]_i_1__0_n_0 ,\current_count_reg[32]_i_1__0_n_1 ,\current_count_reg[32]_i_1__0_n_2 ,\current_count_reg[32]_i_1__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[32]_i_1__0_n_4 ,\current_count_reg[32]_i_1__0_n_5 ,\current_count_reg[32]_i_1__0_n_6 ,\current_count_reg[32]_i_1__0_n_7 }),
        .S(data14[3:0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[32]_i_1__1 
       (.CI(\current_count_reg[28]_i_1__1_n_0 ),
        .CO({\current_count_reg[32]_i_1__1_n_0 ,\current_count_reg[32]_i_1__1_n_1 ,\current_count_reg[32]_i_1__1_n_2 ,\current_count_reg[32]_i_1__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[32]_i_1__1_n_4 ,\current_count_reg[32]_i_1__1_n_5 ,\current_count_reg[32]_i_1__1_n_6 ,\current_count_reg[32]_i_1__1_n_7 }),
        .S(data16[3:0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[36]_i_1 
       (.CI(\current_count_reg[32]_i_1_n_0 ),
        .CO({\current_count_reg[36]_i_1_n_0 ,\current_count_reg[36]_i_1_n_1 ,\current_count_reg[36]_i_1_n_2 ,\current_count_reg[36]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[36]_i_1_n_4 ,\current_count_reg[36]_i_1_n_5 ,\current_count_reg[36]_i_1_n_6 ,\current_count_reg[36]_i_1_n_7 }),
        .S(data12[7:4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[36]_i_1__0 
       (.CI(\current_count_reg[32]_i_1__0_n_0 ),
        .CO({\current_count_reg[36]_i_1__0_n_0 ,\current_count_reg[36]_i_1__0_n_1 ,\current_count_reg[36]_i_1__0_n_2 ,\current_count_reg[36]_i_1__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[36]_i_1__0_n_4 ,\current_count_reg[36]_i_1__0_n_5 ,\current_count_reg[36]_i_1__0_n_6 ,\current_count_reg[36]_i_1__0_n_7 }),
        .S(data14[7:4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[36]_i_1__1 
       (.CI(\current_count_reg[32]_i_1__1_n_0 ),
        .CO({\current_count_reg[36]_i_1__1_n_0 ,\current_count_reg[36]_i_1__1_n_1 ,\current_count_reg[36]_i_1__1_n_2 ,\current_count_reg[36]_i_1__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[36]_i_1__1_n_4 ,\current_count_reg[36]_i_1__1_n_5 ,\current_count_reg[36]_i_1__1_n_6 ,\current_count_reg[36]_i_1__1_n_7 }),
        .S(data16[7:4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[40]_i_1 
       (.CI(\current_count_reg[36]_i_1_n_0 ),
        .CO({\current_count_reg[40]_i_1_n_0 ,\current_count_reg[40]_i_1_n_1 ,\current_count_reg[40]_i_1_n_2 ,\current_count_reg[40]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[40]_i_1_n_4 ,\current_count_reg[40]_i_1_n_5 ,\current_count_reg[40]_i_1_n_6 ,\current_count_reg[40]_i_1_n_7 }),
        .S(data12[11:8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[40]_i_1__0 
       (.CI(\current_count_reg[36]_i_1__0_n_0 ),
        .CO({\current_count_reg[40]_i_1__0_n_0 ,\current_count_reg[40]_i_1__0_n_1 ,\current_count_reg[40]_i_1__0_n_2 ,\current_count_reg[40]_i_1__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[40]_i_1__0_n_4 ,\current_count_reg[40]_i_1__0_n_5 ,\current_count_reg[40]_i_1__0_n_6 ,\current_count_reg[40]_i_1__0_n_7 }),
        .S(data14[11:8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[40]_i_1__1 
       (.CI(\current_count_reg[36]_i_1__1_n_0 ),
        .CO({\current_count_reg[40]_i_1__1_n_0 ,\current_count_reg[40]_i_1__1_n_1 ,\current_count_reg[40]_i_1__1_n_2 ,\current_count_reg[40]_i_1__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[40]_i_1__1_n_4 ,\current_count_reg[40]_i_1__1_n_5 ,\current_count_reg[40]_i_1__1_n_6 ,\current_count_reg[40]_i_1__1_n_7 }),
        .S(data16[11:8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[44]_i_1 
       (.CI(\current_count_reg[40]_i_1_n_0 ),
        .CO({\current_count_reg[44]_i_1_n_0 ,\current_count_reg[44]_i_1_n_1 ,\current_count_reg[44]_i_1_n_2 ,\current_count_reg[44]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[44]_i_1_n_4 ,\current_count_reg[44]_i_1_n_5 ,\current_count_reg[44]_i_1_n_6 ,\current_count_reg[44]_i_1_n_7 }),
        .S(data12[15:12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[44]_i_1__0 
       (.CI(\current_count_reg[40]_i_1__0_n_0 ),
        .CO({\current_count_reg[44]_i_1__0_n_0 ,\current_count_reg[44]_i_1__0_n_1 ,\current_count_reg[44]_i_1__0_n_2 ,\current_count_reg[44]_i_1__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[44]_i_1__0_n_4 ,\current_count_reg[44]_i_1__0_n_5 ,\current_count_reg[44]_i_1__0_n_6 ,\current_count_reg[44]_i_1__0_n_7 }),
        .S(data14[15:12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[44]_i_1__1 
       (.CI(\current_count_reg[40]_i_1__1_n_0 ),
        .CO({\current_count_reg[44]_i_1__1_n_0 ,\current_count_reg[44]_i_1__1_n_1 ,\current_count_reg[44]_i_1__1_n_2 ,\current_count_reg[44]_i_1__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[44]_i_1__1_n_4 ,\current_count_reg[44]_i_1__1_n_5 ,\current_count_reg[44]_i_1__1_n_6 ,\current_count_reg[44]_i_1__1_n_7 }),
        .S(data16[15:12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[48]_i_1 
       (.CI(\current_count_reg[44]_i_1_n_0 ),
        .CO({\current_count_reg[48]_i_1_n_0 ,\current_count_reg[48]_i_1_n_1 ,\current_count_reg[48]_i_1_n_2 ,\current_count_reg[48]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[48]_i_1_n_4 ,\current_count_reg[48]_i_1_n_5 ,\current_count_reg[48]_i_1_n_6 ,\current_count_reg[48]_i_1_n_7 }),
        .S(data12[19:16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[48]_i_1__0 
       (.CI(\current_count_reg[44]_i_1__0_n_0 ),
        .CO({\current_count_reg[48]_i_1__0_n_0 ,\current_count_reg[48]_i_1__0_n_1 ,\current_count_reg[48]_i_1__0_n_2 ,\current_count_reg[48]_i_1__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[48]_i_1__0_n_4 ,\current_count_reg[48]_i_1__0_n_5 ,\current_count_reg[48]_i_1__0_n_6 ,\current_count_reg[48]_i_1__0_n_7 }),
        .S(data14[19:16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[48]_i_1__1 
       (.CI(\current_count_reg[44]_i_1__1_n_0 ),
        .CO({\current_count_reg[48]_i_1__1_n_0 ,\current_count_reg[48]_i_1__1_n_1 ,\current_count_reg[48]_i_1__1_n_2 ,\current_count_reg[48]_i_1__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[48]_i_1__1_n_4 ,\current_count_reg[48]_i_1__1_n_5 ,\current_count_reg[48]_i_1__1_n_6 ,\current_count_reg[48]_i_1__1_n_7 }),
        .S(data16[19:16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[4]_i_1 
       (.CI(\current_count_reg[0]_i_1_n_0 ),
        .CO({\current_count_reg[4]_i_1_n_0 ,\current_count_reg[4]_i_1_n_1 ,\current_count_reg[4]_i_1_n_2 ,\current_count_reg[4]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[4]_i_1_n_4 ,\current_count_reg[4]_i_1_n_5 ,\current_count_reg[4]_i_1_n_6 ,\current_count_reg[4]_i_1_n_7 }),
        .S({\processor/csr_unit/timer_counter/current_count_reg_n_0_[7] ,\processor/csr_unit/timer_counter/current_count_reg_n_0_[6] ,\processor/csr_unit/timer_counter/current_count_reg_n_0_[5] ,\processor/csr_unit/timer_counter/current_count_reg_n_0_[4] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[4]_i_1__0 
       (.CI(current_count_reg[3]),
        .CO({\current_count_reg[4]_i_1__0_n_0 ,\current_count_reg[4]_i_1__0_n_1 ,\current_count_reg[4]_i_1__0_n_2 ,\current_count_reg[4]_i_1__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[4]_i_1__0_n_4 ,\current_count_reg[4]_i_1__0_n_5 ,\current_count_reg[4]_i_1__0_n_6 ,\current_count_reg[4]_i_1__0_n_7 }),
        .S({\processor/csr_unit/cycle_counter/current_count_reg_n_0_[7] ,\processor/csr_unit/cycle_counter/current_count_reg_n_0_[6] ,\processor/csr_unit/cycle_counter/current_count_reg_n_0_[5] ,\processor/csr_unit/cycle_counter/current_count_reg_n_0_[4] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[4]_i_1__1 
       (.CI(\current_count_reg[0]_i_1__1_n_0 ),
        .CO({\current_count_reg[4]_i_1__1_n_0 ,\current_count_reg[4]_i_1__1_n_1 ,\current_count_reg[4]_i_1__1_n_2 ,\current_count_reg[4]_i_1__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[4]_i_1__1_n_4 ,\current_count_reg[4]_i_1__1_n_5 ,\current_count_reg[4]_i_1__1_n_6 ,\current_count_reg[4]_i_1__1_n_7 }),
        .S({\processor/csr_unit/instret_counter/current_count_reg_n_0_[7] ,\processor/csr_unit/instret_counter/current_count_reg_n_0_[6] ,\processor/csr_unit/instret_counter/current_count_reg_n_0_[5] ,\processor/csr_unit/instret_counter/current_count_reg_n_0_[4] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[52]_i_1 
       (.CI(\current_count_reg[48]_i_1_n_0 ),
        .CO({\current_count_reg[52]_i_1_n_0 ,\current_count_reg[52]_i_1_n_1 ,\current_count_reg[52]_i_1_n_2 ,\current_count_reg[52]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[52]_i_1_n_4 ,\current_count_reg[52]_i_1_n_5 ,\current_count_reg[52]_i_1_n_6 ,\current_count_reg[52]_i_1_n_7 }),
        .S(data12[23:20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[52]_i_1__0 
       (.CI(\current_count_reg[48]_i_1__0_n_0 ),
        .CO({\current_count_reg[52]_i_1__0_n_0 ,\current_count_reg[52]_i_1__0_n_1 ,\current_count_reg[52]_i_1__0_n_2 ,\current_count_reg[52]_i_1__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[52]_i_1__0_n_4 ,\current_count_reg[52]_i_1__0_n_5 ,\current_count_reg[52]_i_1__0_n_6 ,\current_count_reg[52]_i_1__0_n_7 }),
        .S(data14[23:20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[52]_i_1__1 
       (.CI(\current_count_reg[48]_i_1__1_n_0 ),
        .CO({\current_count_reg[52]_i_1__1_n_0 ,\current_count_reg[52]_i_1__1_n_1 ,\current_count_reg[52]_i_1__1_n_2 ,\current_count_reg[52]_i_1__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[52]_i_1__1_n_4 ,\current_count_reg[52]_i_1__1_n_5 ,\current_count_reg[52]_i_1__1_n_6 ,\current_count_reg[52]_i_1__1_n_7 }),
        .S(data16[23:20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[56]_i_1 
       (.CI(\current_count_reg[52]_i_1_n_0 ),
        .CO({\current_count_reg[56]_i_1_n_0 ,\current_count_reg[56]_i_1_n_1 ,\current_count_reg[56]_i_1_n_2 ,\current_count_reg[56]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[56]_i_1_n_4 ,\current_count_reg[56]_i_1_n_5 ,\current_count_reg[56]_i_1_n_6 ,\current_count_reg[56]_i_1_n_7 }),
        .S(data12[27:24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[56]_i_1__0 
       (.CI(\current_count_reg[52]_i_1__0_n_0 ),
        .CO({\current_count_reg[56]_i_1__0_n_0 ,\current_count_reg[56]_i_1__0_n_1 ,\current_count_reg[56]_i_1__0_n_2 ,\current_count_reg[56]_i_1__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[56]_i_1__0_n_4 ,\current_count_reg[56]_i_1__0_n_5 ,\current_count_reg[56]_i_1__0_n_6 ,\current_count_reg[56]_i_1__0_n_7 }),
        .S(data14[27:24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[56]_i_1__1 
       (.CI(\current_count_reg[52]_i_1__1_n_0 ),
        .CO({\current_count_reg[56]_i_1__1_n_0 ,\current_count_reg[56]_i_1__1_n_1 ,\current_count_reg[56]_i_1__1_n_2 ,\current_count_reg[56]_i_1__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[56]_i_1__1_n_4 ,\current_count_reg[56]_i_1__1_n_5 ,\current_count_reg[56]_i_1__1_n_6 ,\current_count_reg[56]_i_1__1_n_7 }),
        .S(data16[27:24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[60]_i_1 
       (.CI(\current_count_reg[56]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[60]_i_1_n_4 ,\current_count_reg[60]_i_1_n_5 ,\current_count_reg[60]_i_1_n_6 ,\current_count_reg[60]_i_1_n_7 }),
        .S(data12[31:28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[60]_i_1__0 
       (.CI(\current_count_reg[56]_i_1__0_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[60]_i_1__0_n_4 ,\current_count_reg[60]_i_1__0_n_5 ,\current_count_reg[60]_i_1__0_n_6 ,\current_count_reg[60]_i_1__0_n_7 }),
        .S(data14[31:28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[60]_i_1__1 
       (.CI(\current_count_reg[56]_i_1__1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[60]_i_1__1_n_4 ,\current_count_reg[60]_i_1__1_n_5 ,\current_count_reg[60]_i_1__1_n_6 ,\current_count_reg[60]_i_1__1_n_7 }),
        .S(data16[31:28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[8]_i_1 
       (.CI(\current_count_reg[4]_i_1_n_0 ),
        .CO({\current_count_reg[8]_i_1_n_0 ,\current_count_reg[8]_i_1_n_1 ,\current_count_reg[8]_i_1_n_2 ,\current_count_reg[8]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[8]_i_1_n_4 ,\current_count_reg[8]_i_1_n_5 ,\current_count_reg[8]_i_1_n_6 ,\current_count_reg[8]_i_1_n_7 }),
        .S({\processor/csr_unit/timer_counter/current_count_reg_n_0_[11] ,\processor/csr_unit/timer_counter/current_count_reg_n_0_[10] ,\processor/csr_unit/timer_counter/current_count_reg_n_0_[9] ,\processor/csr_unit/timer_counter/current_count_reg_n_0_[8] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[8]_i_1__0 
       (.CI(\current_count_reg[4]_i_1__0_n_0 ),
        .CO({\current_count_reg[8]_i_1__0_n_0 ,\current_count_reg[8]_i_1__0_n_1 ,\current_count_reg[8]_i_1__0_n_2 ,\current_count_reg[8]_i_1__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[8]_i_1__0_n_4 ,\current_count_reg[8]_i_1__0_n_5 ,\current_count_reg[8]_i_1__0_n_6 ,\current_count_reg[8]_i_1__0_n_7 }),
        .S({\processor/csr_unit/cycle_counter/current_count_reg_n_0_[11] ,\processor/csr_unit/cycle_counter/current_count_reg_n_0_[10] ,\processor/csr_unit/cycle_counter/current_count_reg_n_0_[9] ,\processor/csr_unit/cycle_counter/current_count_reg_n_0_[8] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \current_count_reg[8]_i_1__1 
       (.CI(\current_count_reg[4]_i_1__1_n_0 ),
        .CO({\current_count_reg[8]_i_1__1_n_0 ,\current_count_reg[8]_i_1__1_n_1 ,\current_count_reg[8]_i_1__1_n_2 ,\current_count_reg[8]_i_1__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\current_count_reg[8]_i_1__1_n_4 ,\current_count_reg[8]_i_1__1_n_5 ,\current_count_reg[8]_i_1__1_n_6 ,\current_count_reg[8]_i_1__1_n_7 }),
        .S({\processor/csr_unit/instret_counter/current_count_reg_n_0_[11] ,\processor/csr_unit/instret_counter/current_count_reg_n_0_[10] ,\processor/csr_unit/instret_counter/current_count_reg_n_0_[9] ,\processor/csr_unit/instret_counter/current_count_reg_n_0_[8] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A0A2AA00000200)) 
    \decode_exception_cause[0]_i_1 
       (.I0(decode_exception_cause),
        .I1(\processor/decode/instruction_reg_n_0_[3] ),
        .I2(\decode_exception_cause[0]_i_3_n_0 ),
        .I3(\processor/decode/instruction_reg_n_0_[4] ),
        .I4(\processor/decode/instruction_reg_n_0_[6] ),
        .I5(\decode_exception_cause[3]_i_4_n_0 ),
        .O(\processor/id_exception_cause [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAA8AAAA)) 
    \decode_exception_cause[0]_i_2 
       (.I0(decode_exception_cause1),
        .I1(\branch[2]_i_4_n_0 ),
        .I2(\processor/id_shamt [1]),
        .I3(\processor/id_csr_use_immediate ),
        .I4(\decode_exception_cause[0]_i_4_n_0 ),
        .I5(\decode_exception_cause[0]_i_5_n_0 ),
        .O(decode_exception_cause));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF01000000000000)) 
    \decode_exception_cause[0]_i_3 
       (.I0(data0[31]),
        .I1(data0[30]),
        .I2(\decode_exception_cause[0]_i_6_n_0 ),
        .I3(\decode_exception_cause[3]_i_5_n_0 ),
        .I4(\processor/decode/instruction_reg_n_0_[6] ),
        .I5(\processor/decode/instruction_reg_n_0_[5] ),
        .O(\decode_exception_cause[0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \decode_exception_cause[0]_i_4 
       (.I0(\processor/id_shamt [3]),
        .I1(\processor/id_shamt [2]),
        .O(\decode_exception_cause[0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF7FFF)) 
    \decode_exception_cause[0]_i_5 
       (.I0(\processor/decode/instruction_reg_n_0_[6] ),
        .I1(data0[28]),
        .I2(\processor/decode/instruction_reg_n_0_[4] ),
        .I3(\processor/id_shamt [0]),
        .I4(\processor/decode/instruction_reg_n_0_ ),
        .I5(\decode_exception_cause[0]_i_7_n_0 ),
        .O(\decode_exception_cause[0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \decode_exception_cause[0]_i_6 
       (.I0(data0[26]),
        .I1(data0[25]),
        .I2(data0[29]),
        .I3(data0[27]),
        .I4(\decode_exception_cause[0]_i_8_n_0 ),
        .O(\decode_exception_cause[0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \decode_exception_cause[0]_i_7 
       (.I0(\processor/id_funct3 [1]),
        .I1(\processor/id_funct3 [0]),
        .O(\decode_exception_cause[0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \decode_exception_cause[0]_i_8 
       (.I0(\processor/id_shamt [3]),
        .I1(\processor/id_shamt [4]),
        .I2(\processor/id_shamt [1]),
        .I3(\processor/id_shamt [2]),
        .O(\decode_exception_cause[0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAA22A200002202)) 
    \decode_exception_cause[2]_i_1 
       (.I0(decode_exception_cause1),
        .I1(\immediate[30]_i_2_n_0 ),
        .I2(\decode_exception_cause[2]_i_2_n_0 ),
        .I3(\decode_exception_cause[2]_i_3_n_0 ),
        .I4(\decode_exception_cause[2]_i_4_n_0 ),
        .I5(\decode_exception_cause[3]_i_4_n_0 ),
        .O(\processor/id_exception_cause [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAAB)) 
    \decode_exception_cause[2]_i_2 
       (.I0(\decode_exception_cause[3]_i_5_n_0 ),
        .I1(\decode_exception_cause[2]_i_5_n_0 ),
        .I2(data0[31]),
        .I3(data0[30]),
        .I4(\processor/id_shamt [0]),
        .I5(data0[29]),
        .O(\decode_exception_cause[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \decode_exception_cause[2]_i_3 
       (.I0(\processor/decode/instruction_reg_n_0_[5] ),
        .I1(\processor/decode/instruction_reg_n_0_[6] ),
        .O(\decode_exception_cause[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \decode_exception_cause[2]_i_4 
       (.I0(\processor/decode/instruction_reg_n_0_[4] ),
        .I1(\processor/decode/instruction_reg_n_0_[6] ),
        .O(\decode_exception_cause[2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFEFFFF)) 
    \decode_exception_cause[2]_i_5 
       (.I0(\branch[2]_i_4_n_0 ),
        .I1(\processor/id_shamt [3]),
        .I2(\processor/id_shamt [2]),
        .I3(\processor/id_shamt [1]),
        .I4(data0[28]),
        .O(\decode_exception_cause[2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A0A2AA00000200)) 
    \decode_exception_cause[3]_i_1 
       (.I0(decode_exception_cause1),
        .I1(\processor/decode/instruction_reg_n_0_[3] ),
        .I2(\decode_exception_cause[3]_i_3_n_0 ),
        .I3(\processor/decode/instruction_reg_n_0_[4] ),
        .I4(\processor/decode/instruction_reg_n_0_[6] ),
        .I5(\decode_exception_cause[3]_i_4_n_0 ),
        .O(\processor/id_exception_cause [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF7)) 
    \decode_exception_cause[3]_i_2 
       (.I0(\processor/id_alu_op [1]),
        .I1(\processor/id_alu_op [0]),
        .I2(decode_exception_i_5_n_0),
        .O(decode_exception_cause1));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFF0001)) 
    \decode_exception_cause[3]_i_3 
       (.I0(data0[31]),
        .I1(data0[29]),
        .I2(data0[30]),
        .I3(decode_exception_i_4_n_0),
        .I4(\decode_exception_cause[3]_i_5_n_0 ),
        .I5(\decode_exception_cause[2]_i_3_n_0 ),
        .O(\decode_exception_cause[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h220FF20F)) 
    \decode_exception_cause[3]_i_4 
       (.I0(\processor/decode/instruction_reg_n_0_[6] ),
        .I1(\processor/decode/instruction_reg_n_0_[4] ),
        .I2(\processor/decode/instruction_reg_n_0_[3] ),
        .I3(\processor/decode/instruction_reg_n_0_ ),
        .I4(\processor/decode/instruction_reg_n_0_[5] ),
        .O(\decode_exception_cause[3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFD)) 
    \decode_exception_cause[3]_i_5 
       (.I0(\processor/decode/instruction_reg_n_0_[4] ),
        .I1(\processor/id_csr_use_immediate ),
        .I2(\processor/id_funct3 [0]),
        .I3(\processor/id_funct3 [1]),
        .O(\decode_exception_cause[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA8A8A8A8FFA8A8A8)) 
    decode_exception_i_1
       (.I0(decode_exception_i_2_n_0),
        .I1(decode_exception_i_3_n_0),
        .I2(decode_exception_i_4_n_0),
        .I3(\processor/id_alu_op [1]),
        .I4(\processor/id_alu_op [0]),
        .I5(decode_exception_i_5_n_0),
        .O(\processor/id_exception ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFCCE6CC44CCE6)) 
    decode_exception_i_2
       (.I0(\processor/decode/instruction_reg_n_0_ ),
        .I1(\processor/decode/instruction_reg_n_0_[3] ),
        .I2(\processor/decode/instruction_reg_n_0_[5] ),
        .I3(\processor/decode/instruction_reg_n_0_[4] ),
        .I4(\processor/decode/instruction_reg_n_0_[6] ),
        .I5(decode_exception_i_6_n_0),
        .O(decode_exception_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFDF)) 
    decode_exception_i_3
       (.I0(\processor/decode/instruction_reg_n_0_[5] ),
        .I1(\processor/decode/instruction_reg_n_0_[3] ),
        .I2(data0[28]),
        .I3(data0[29]),
        .I4(\processor/decode/instruction_reg_n_0_ ),
        .I5(decode_exception_i_7_n_0),
        .O(decode_exception_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    decode_exception_i_4
       (.I0(\branch[2]_i_4_n_0 ),
        .I1(\processor/id_shamt [1]),
        .I2(\processor/id_shamt [0]),
        .I3(\processor/id_shamt [3]),
        .I4(\processor/id_shamt [2]),
        .O(decode_exception_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    decode_exception_i_5
       (.I0(\processor/id_alu_op [2]),
        .I1(\processor/id_alu_op [3]),
        .O(decode_exception_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDDDDDDF55555555)) 
    decode_exception_i_6
       (.I0(\processor/decode/instruction_reg_n_0_[5] ),
        .I1(\processor/decode/instruction_reg_n_0_ ),
        .I2(\processor/id_csr_use_immediate ),
        .I3(\processor/id_funct3 [0]),
        .I4(\processor/id_funct3 [1]),
        .I5(\processor/decode/instruction_reg_n_0_[4] ),
        .O(decode_exception_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    decode_exception_i_7
       (.I0(data0[31]),
        .I1(data0[30]),
        .O(decode_exception_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \dmem_address_p[31]_i_1 
       (.I0(\dmem_address_p[31]_i_2_n_0 ),
        .I1(\processor/memory/p_1_in ),
        .O(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF1)) 
    \dmem_address_p[31]_i_2 
       (.I0(\processor/ex_mem_op [1]),
        .I1(\processor/ex_mem_op [2]),
        .I2(\mem_op[2]_i_5_n_0 ),
        .O(\dmem_address_p[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair148" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \dmem_data_out[0]_i_1 
       (.I0(\dmem_data_out[8]_i_2_n_0 ),
        .I1(\dmem_data_out[23]_i_3_n_0 ),
        .I2(dmem_data_out),
        .O(SHIFT_RIGHT[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000B080)) 
    \dmem_data_out[0]_i_2 
       (.I0(wb_dat_in[16]),
        .I1(\dmem_data_out[23]_i_4_n_0 ),
        .I2(\arbiter/state [1]),
        .I3(wb_dat_in[0]),
        .I4(\arbiter/state [0]),
        .O(dmem_data_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0040FFFF00400000)) 
    \dmem_data_out[10]_i_1 
       (.I0(\arbiter/state [0]),
        .I1(wb_dat_in[18]),
        .I2(\arbiter/state [1]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .I4(\dmem_data_out[23]_i_3_n_0 ),
        .I5(\dmem_data_out[10]_i_2_n_0 ),
        .O(SHIFT_RIGHT[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000B080)) 
    \dmem_data_out[10]_i_2 
       (.I0(wb_dat_in[26]),
        .I1(\dmem_data_out[23]_i_4_n_0 ),
        .I2(\arbiter/state [1]),
        .I3(wb_dat_in[10]),
        .I4(\arbiter/state [0]),
        .O(\dmem_data_out[10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0040FFFF00400000)) 
    \dmem_data_out[11]_i_1 
       (.I0(\arbiter/state [0]),
        .I1(wb_dat_in[19]),
        .I2(\arbiter/state [1]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .I4(\dmem_data_out[23]_i_3_n_0 ),
        .I5(\dmem_data_out[11]_i_2_n_0 ),
        .O(SHIFT_RIGHT[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000B080)) 
    \dmem_data_out[11]_i_2 
       (.I0(wb_dat_in[27]),
        .I1(\dmem_data_out[23]_i_4_n_0 ),
        .I2(\arbiter/state [1]),
        .I3(wb_dat_in[11]),
        .I4(\arbiter/state [0]),
        .O(\dmem_data_out[11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0040FFFF00400000)) 
    \dmem_data_out[12]_i_1 
       (.I0(\arbiter/state [0]),
        .I1(wb_dat_in[20]),
        .I2(\arbiter/state [1]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .I4(\dmem_data_out[23]_i_3_n_0 ),
        .I5(\dmem_data_out[12]_i_2_n_0 ),
        .O(SHIFT_RIGHT[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000B080)) 
    \dmem_data_out[12]_i_2 
       (.I0(wb_dat_in[28]),
        .I1(\dmem_data_out[23]_i_4_n_0 ),
        .I2(\arbiter/state [1]),
        .I3(wb_dat_in[12]),
        .I4(\arbiter/state [0]),
        .O(\dmem_data_out[12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0040FFFF00400000)) 
    \dmem_data_out[13]_i_1 
       (.I0(\arbiter/state [0]),
        .I1(wb_dat_in[21]),
        .I2(\arbiter/state [1]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .I4(\dmem_data_out[23]_i_3_n_0 ),
        .I5(\dmem_data_out[13]_i_2_n_0 ),
        .O(SHIFT_RIGHT[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000B080)) 
    \dmem_data_out[13]_i_2 
       (.I0(wb_dat_in[29]),
        .I1(\dmem_data_out[23]_i_4_n_0 ),
        .I2(\arbiter/state [1]),
        .I3(wb_dat_in[13]),
        .I4(\arbiter/state [0]),
        .O(\dmem_data_out[13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0040FFFF00400000)) 
    \dmem_data_out[14]_i_1 
       (.I0(\arbiter/state [0]),
        .I1(wb_dat_in[22]),
        .I2(\arbiter/state [1]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .I4(\dmem_data_out[23]_i_3_n_0 ),
        .I5(\dmem_data_out[14]_i_2_n_0 ),
        .O(SHIFT_RIGHT[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000B080)) 
    \dmem_data_out[14]_i_2 
       (.I0(wb_dat_in[30]),
        .I1(\dmem_data_out[23]_i_4_n_0 ),
        .I2(\arbiter/state [1]),
        .I3(wb_dat_in[14]),
        .I4(\arbiter/state [0]),
        .O(\dmem_data_out[14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0040FFFF00400000)) 
    \dmem_data_out[15]_i_1 
       (.I0(\arbiter/state [0]),
        .I1(wb_dat_in[23]),
        .I2(\arbiter/state [1]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .I4(\dmem_data_out[23]_i_3_n_0 ),
        .I5(\dmem_data_out[15]_i_2_n_0 ),
        .O(SHIFT_RIGHT[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000B080)) 
    \dmem_data_out[15]_i_2 
       (.I0(wb_dat_in[31]),
        .I1(\dmem_data_out[23]_i_4_n_0 ),
        .I2(\arbiter/state [1]),
        .I3(wb_dat_in[15]),
        .I4(\arbiter/state [0]),
        .O(\dmem_data_out[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000B080000)) 
    \dmem_data_out[16]_i_1 
       (.I0(wb_dat_in[24]),
        .I1(\dmem_data_out[23]_i_3_n_0 ),
        .I2(\arbiter/state [0]),
        .I3(wb_dat_in[16]),
        .I4(\arbiter/state [1]),
        .I5(\dmem_data_out[23]_i_4_n_0 ),
        .O(SHIFT_RIGHT[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000B080000)) 
    \dmem_data_out[17]_i_1 
       (.I0(wb_dat_in[25]),
        .I1(\dmem_data_out[23]_i_3_n_0 ),
        .I2(\arbiter/state [0]),
        .I3(wb_dat_in[17]),
        .I4(\arbiter/state [1]),
        .I5(\dmem_data_out[23]_i_4_n_0 ),
        .O(SHIFT_RIGHT[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000B080000)) 
    \dmem_data_out[18]_i_1 
       (.I0(wb_dat_in[26]),
        .I1(\dmem_data_out[23]_i_3_n_0 ),
        .I2(\arbiter/state [0]),
        .I3(wb_dat_in[18]),
        .I4(\arbiter/state [1]),
        .I5(\dmem_data_out[23]_i_4_n_0 ),
        .O(SHIFT_RIGHT[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000B080000)) 
    \dmem_data_out[19]_i_1 
       (.I0(wb_dat_in[27]),
        .I1(\dmem_data_out[23]_i_3_n_0 ),
        .I2(\arbiter/state [0]),
        .I3(wb_dat_in[19]),
        .I4(\arbiter/state [1]),
        .I5(\dmem_data_out[23]_i_4_n_0 ),
        .O(SHIFT_RIGHT[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair148" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \dmem_data_out[1]_i_1 
       (.I0(\dmem_data_out[9]_i_2_n_0 ),
        .I1(\dmem_data_out[23]_i_3_n_0 ),
        .I2(\dmem_data_out[1]_i_2_n_0 ),
        .O(SHIFT_RIGHT[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000B080)) 
    \dmem_data_out[1]_i_2 
       (.I0(wb_dat_in[17]),
        .I1(\dmem_data_out[23]_i_4_n_0 ),
        .I2(\arbiter/state [1]),
        .I3(wb_dat_in[1]),
        .I4(\arbiter/state [0]),
        .O(\dmem_data_out[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000B080000)) 
    \dmem_data_out[20]_i_1 
       (.I0(wb_dat_in[28]),
        .I1(\dmem_data_out[23]_i_3_n_0 ),
        .I2(\arbiter/state [0]),
        .I3(wb_dat_in[20]),
        .I4(\arbiter/state [1]),
        .I5(\dmem_data_out[23]_i_4_n_0 ),
        .O(SHIFT_RIGHT[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000B080000)) 
    \dmem_data_out[21]_i_1 
       (.I0(wb_dat_in[29]),
        .I1(\dmem_data_out[23]_i_3_n_0 ),
        .I2(\arbiter/state [0]),
        .I3(wb_dat_in[21]),
        .I4(\arbiter/state [1]),
        .I5(\dmem_data_out[23]_i_4_n_0 ),
        .O(SHIFT_RIGHT[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000B080000)) 
    \dmem_data_out[22]_i_1 
       (.I0(wb_dat_in[30]),
        .I1(\dmem_data_out[23]_i_3_n_0 ),
        .I2(\arbiter/state [0]),
        .I3(wb_dat_in[22]),
        .I4(\arbiter/state [1]),
        .I5(\dmem_data_out[23]_i_4_n_0 ),
        .O(SHIFT_RIGHT[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00004000)) 
    \dmem_data_out[23]_i_1 
       (.I0(\arbiter/state [0]),
        .I1(wb_ack_in),
        .I2(\arbiter/state [1]),
        .I3(\dmem_if/state_reg_n_0_ ),
        .I4(reset),
        .O(\dmem_data_out[23]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000B080000)) 
    \dmem_data_out[23]_i_2 
       (.I0(wb_dat_in[31]),
        .I1(\dmem_data_out[23]_i_3_n_0 ),
        .I2(\arbiter/state [0]),
        .I3(wb_dat_in[23]),
        .I4(\arbiter/state [1]),
        .I5(\dmem_data_out[23]_i_4_n_0 ),
        .O(SHIFT_RIGHT[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h004000400040CC40)) 
    \dmem_data_out[23]_i_3 
       (.I0(\processor/dmem_data_size_p [1]),
        .I1(dmem_address[0]),
        .I2(\processor/dmem_data_size_p [0]),
        .I3(\processor/memory/p_1_in ),
        .I4(\processor/ex_dmem_data_size [1]),
        .I5(\processor/ex_mem_size ),
        .O(\dmem_data_out[23]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h75200000)) 
    \dmem_data_out[23]_i_4 
       (.I0(\processor/memory/p_1_in ),
        .I1(\dmem_address_p[31]_i_2_n_0 ),
        .I2(\processor/ex_rd_data [1]),
        .I3(dmem_address_p[1]),
        .I4(\dmem_data_out[23]_i_5_n_0 ),
        .O(\dmem_data_out[23]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h535C)) 
    \dmem_data_out[23]_i_5 
       (.I0(\processor/ex_mem_size ),
        .I1(\processor/dmem_data_size_p [0]),
        .I2(\processor/memory/p_1_in ),
        .I3(\processor/dmem_data_size_p [1]),
        .O(\dmem_data_out[23]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \dmem_data_out[24]_i_1 
       (.I0(\arbiter/state [0]),
        .I1(wb_dat_in[24]),
        .I2(\arbiter/state [1]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .O(\dmem_data_out[24]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \dmem_data_out[25]_i_1 
       (.I0(\arbiter/state [0]),
        .I1(wb_dat_in[25]),
        .I2(\arbiter/state [1]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .O(\dmem_data_out[25]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \dmem_data_out[26]_i_1 
       (.I0(\arbiter/state [0]),
        .I1(wb_dat_in[26]),
        .I2(\arbiter/state [1]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .O(\dmem_data_out[26]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \dmem_data_out[27]_i_1 
       (.I0(\arbiter/state [0]),
        .I1(wb_dat_in[27]),
        .I2(\arbiter/state [1]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .O(\dmem_data_out[27]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \dmem_data_out[28]_i_1 
       (.I0(\arbiter/state [0]),
        .I1(wb_dat_in[28]),
        .I2(\arbiter/state [1]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .O(\dmem_data_out[28]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \dmem_data_out[29]_i_1 
       (.I0(\arbiter/state [0]),
        .I1(wb_dat_in[29]),
        .I2(\arbiter/state [1]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .O(\dmem_data_out[29]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair150" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \dmem_data_out[2]_i_1 
       (.I0(\dmem_data_out[10]_i_2_n_0 ),
        .I1(\dmem_data_out[23]_i_3_n_0 ),
        .I2(\dmem_data_out[2]_i_2_n_0 ),
        .O(SHIFT_RIGHT[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000B080)) 
    \dmem_data_out[2]_i_2 
       (.I0(wb_dat_in[18]),
        .I1(\dmem_data_out[23]_i_4_n_0 ),
        .I2(\arbiter/state [1]),
        .I3(wb_dat_in[2]),
        .I4(\arbiter/state [0]),
        .O(\dmem_data_out[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \dmem_data_out[30]_i_1 
       (.I0(\arbiter/state [0]),
        .I1(wb_dat_in[30]),
        .I2(\arbiter/state [1]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .O(\dmem_data_out[30]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \dmem_data_out[31]_i_2 
       (.I0(\arbiter/state [0]),
        .I1(wb_dat_in[31]),
        .I2(\arbiter/state [1]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .O(\dmem_data_out[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair150" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \dmem_data_out[3]_i_1 
       (.I0(\dmem_data_out[11]_i_2_n_0 ),
        .I1(\dmem_data_out[23]_i_3_n_0 ),
        .I2(\dmem_data_out[3]_i_2_n_0 ),
        .O(SHIFT_RIGHT[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000B080)) 
    \dmem_data_out[3]_i_2 
       (.I0(wb_dat_in[19]),
        .I1(\dmem_data_out[23]_i_4_n_0 ),
        .I2(\arbiter/state [1]),
        .I3(wb_dat_in[3]),
        .I4(\arbiter/state [0]),
        .O(\dmem_data_out[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair152" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \dmem_data_out[4]_i_1 
       (.I0(\dmem_data_out[12]_i_2_n_0 ),
        .I1(\dmem_data_out[23]_i_3_n_0 ),
        .I2(\dmem_data_out[4]_i_2_n_0 ),
        .O(SHIFT_RIGHT[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000B080)) 
    \dmem_data_out[4]_i_2 
       (.I0(wb_dat_in[20]),
        .I1(\dmem_data_out[23]_i_4_n_0 ),
        .I2(\arbiter/state [1]),
        .I3(wb_dat_in[4]),
        .I4(\arbiter/state [0]),
        .O(\dmem_data_out[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair152" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \dmem_data_out[5]_i_1 
       (.I0(\dmem_data_out[13]_i_2_n_0 ),
        .I1(\dmem_data_out[23]_i_3_n_0 ),
        .I2(\dmem_data_out[5]_i_2_n_0 ),
        .O(SHIFT_RIGHT[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000B080)) 
    \dmem_data_out[5]_i_2 
       (.I0(wb_dat_in[21]),
        .I1(\dmem_data_out[23]_i_4_n_0 ),
        .I2(\arbiter/state [1]),
        .I3(wb_dat_in[5]),
        .I4(\arbiter/state [0]),
        .O(\dmem_data_out[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \dmem_data_out[6]_i_1 
       (.I0(\dmem_data_out[14]_i_2_n_0 ),
        .I1(\dmem_data_out[23]_i_3_n_0 ),
        .I2(\dmem_data_out[6]_i_2_n_0 ),
        .O(SHIFT_RIGHT[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000B080)) 
    \dmem_data_out[6]_i_2 
       (.I0(wb_dat_in[22]),
        .I1(\dmem_data_out[23]_i_4_n_0 ),
        .I2(\arbiter/state [1]),
        .I3(wb_dat_in[6]),
        .I4(\arbiter/state [0]),
        .O(\dmem_data_out[6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \dmem_data_out[7]_i_1 
       (.I0(\dmem_data_out[15]_i_2_n_0 ),
        .I1(\dmem_data_out[23]_i_3_n_0 ),
        .I2(\dmem_data_out[7]_i_2_n_0 ),
        .O(SHIFT_RIGHT[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000B080)) 
    \dmem_data_out[7]_i_2 
       (.I0(wb_dat_in[23]),
        .I1(\dmem_data_out[23]_i_4_n_0 ),
        .I2(\arbiter/state [1]),
        .I3(wb_dat_in[7]),
        .I4(\arbiter/state [0]),
        .O(\dmem_data_out[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0040FFFF00400000)) 
    \dmem_data_out[8]_i_1 
       (.I0(\arbiter/state [0]),
        .I1(wb_dat_in[16]),
        .I2(\arbiter/state [1]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .I4(\dmem_data_out[23]_i_3_n_0 ),
        .I5(\dmem_data_out[8]_i_2_n_0 ),
        .O(SHIFT_RIGHT[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000B080)) 
    \dmem_data_out[8]_i_2 
       (.I0(wb_dat_in[24]),
        .I1(\dmem_data_out[23]_i_4_n_0 ),
        .I2(\arbiter/state [1]),
        .I3(wb_dat_in[8]),
        .I4(\arbiter/state [0]),
        .O(\dmem_data_out[8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0040FFFF00400000)) 
    \dmem_data_out[9]_i_1 
       (.I0(\arbiter/state [0]),
        .I1(wb_dat_in[17]),
        .I2(\arbiter/state [1]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .I4(\dmem_data_out[23]_i_3_n_0 ),
        .I5(\dmem_data_out[9]_i_2_n_0 ),
        .O(SHIFT_RIGHT[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000B080)) 
    \dmem_data_out[9]_i_2 
       (.I0(wb_dat_in[25]),
        .I1(\dmem_data_out[23]_i_4_n_0 ),
        .I2(\arbiter/state [1]),
        .I3(wb_dat_in[9]),
        .I4(\arbiter/state [0]),
        .O(\dmem_data_out[9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[0]_i_1 
       (.I0(\processor/mem_rd_data [0]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [0]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [0]),
        .O(\processor/ex_dmem_data_out [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[10]_i_1 
       (.I0(\processor/mem_rd_data [10]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [10]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [10]),
        .O(\processor/ex_dmem_data_out [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCAA00AAFFFFFFFF)) 
    \dmem_data_out_p[10]_i_2 
       (.I0(rd_data[10]),
        .I1(\mem_size[0]_repN ),
        .I2(\mem_size[1]_repN ),
        .I3(\rd_data_out[31]_i_4_n_0 ),
        .I4(\dmem_if/dmem_data_out_reg_n_0_[10] ),
        .I5(\rd_data_out[15]_i_3_n_0 ),
        .O(\processor/mem_rd_data [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[11]_i_1 
       (.I0(\processor/mem_rd_data [11]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [11]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [11]),
        .O(\processor/ex_dmem_data_out [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCAA00AAFFFFFFFF)) 
    \dmem_data_out_p[11]_i_2 
       (.I0(rd_data[11]),
        .I1(\mem_size[0]_repN ),
        .I2(\mem_size[1]_repN ),
        .I3(\rd_data_out[31]_i_4_n_0 ),
        .I4(\dmem_if/dmem_data_out_reg_n_0_[11] ),
        .I5(\rd_data_out[15]_i_3_n_0 ),
        .O(\processor/mem_rd_data [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[12]_i_1 
       (.I0(\processor/mem_rd_data [12]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [12]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [12]),
        .O(\processor/ex_dmem_data_out [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCAA00AAFFFFFFFF)) 
    \dmem_data_out_p[12]_i_2 
       (.I0(rd_data[12]),
        .I1(\mem_size[0]_repN ),
        .I2(\mem_size[1]_repN ),
        .I3(\rd_data_out[31]_i_4_n_0 ),
        .I4(\dmem_if/dmem_data_out_reg_n_0_[12] ),
        .I5(\rd_data_out[15]_i_3_n_0 ),
        .O(\processor/mem_rd_data [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[13]_i_1 
       (.I0(\processor/mem_rd_data [13]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [13]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [13]),
        .O(\processor/ex_dmem_data_out [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCAA00AAFFFFFFFF)) 
    \dmem_data_out_p[13]_i_2 
       (.I0(rd_data[13]),
        .I1(\mem_size[0]_repN ),
        .I2(\mem_size[1]_repN ),
        .I3(\rd_data_out[31]_i_4_n_0 ),
        .I4(\dmem_if/dmem_data_out_reg_n_0_[13] ),
        .I5(\rd_data_out[15]_i_3_n_0 ),
        .O(\processor/mem_rd_data [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[14]_i_1 
       (.I0(\processor/mem_rd_data [14]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [14]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [14]),
        .O(\processor/ex_dmem_data_out [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCAA00AAFFFFFFFF)) 
    \dmem_data_out_p[14]_i_2 
       (.I0(rd_data[14]),
        .I1(\mem_size[0]_repN ),
        .I2(\mem_size[1]_repN ),
        .I3(\rd_data_out[31]_i_4_n_0 ),
        .I4(\dmem_if/dmem_data_out_reg_n_0_[14] ),
        .I5(\rd_data_out[15]_i_3_n_0 ),
        .O(\processor/mem_rd_data [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[15]_i_1 
       (.I0(\processor/mem_rd_data [15]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [15]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [15]),
        .O(\processor/ex_dmem_data_out [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCAA00AAFFFFFFFF)) 
    \dmem_data_out_p[15]_i_2 
       (.I0(rd_data[15]),
        .I1(\mem_size[0]_repN ),
        .I2(\mem_size[1]_repN ),
        .I3(\rd_data_out[31]_i_4_n_0 ),
        .I4(p_1_in0),
        .I5(\rd_data_out[15]_i_3_n_0 ),
        .O(\processor/mem_rd_data [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[16]_i_1 
       (.I0(\processor/mem_rd_data [16]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [16]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [16]),
        .O(\processor/ex_dmem_data_out [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[17]_i_1 
       (.I0(\processor/mem_rd_data [17]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [17]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [17]),
        .O(\processor/ex_dmem_data_out [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[18]_i_1 
       (.I0(\processor/mem_rd_data [18]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [18]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [18]),
        .O(\processor/ex_dmem_data_out [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[19]_i_1 
       (.I0(\processor/mem_rd_data [19]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [19]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [19]),
        .O(\processor/ex_dmem_data_out [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[1]_i_1 
       (.I0(\processor/mem_rd_data [1]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [1]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [1]),
        .O(\processor/ex_dmem_data_out [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[20]_i_1 
       (.I0(\processor/mem_rd_data [20]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [20]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [20]),
        .O(\processor/ex_dmem_data_out [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[21]_i_1 
       (.I0(\processor/mem_rd_data [21]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [21]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [21]),
        .O(\processor/ex_dmem_data_out [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[22]_i_1 
       (.I0(\processor/mem_rd_data [22]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [22]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [22]),
        .O(\processor/ex_dmem_data_out [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[23]_i_1 
       (.I0(\processor/mem_rd_data [23]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [23]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [23]),
        .O(\processor/ex_dmem_data_out [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[24]_i_1 
       (.I0(\processor/mem_rd_data [24]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [24]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [24]),
        .O(\processor/ex_dmem_data_out [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[25]_i_1 
       (.I0(\processor/mem_rd_data [25]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [25]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [25]),
        .O(\processor/ex_dmem_data_out [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[26]_i_1 
       (.I0(\processor/mem_rd_data [26]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [26]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [26]),
        .O(\processor/ex_dmem_data_out [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[27]_i_1 
       (.I0(\processor/mem_rd_data [27]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [27]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [27]),
        .O(\processor/ex_dmem_data_out [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[28]_i_1 
       (.I0(\processor/mem_rd_data [28]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [28]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [28]),
        .O(\processor/ex_dmem_data_out [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[29]_i_1 
       (.I0(\processor/mem_rd_data [29]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [29]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [29]),
        .O(\processor/ex_dmem_data_out [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[2]_i_1 
       (.I0(\processor/mem_rd_data [2]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [2]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [2]),
        .O(\processor/ex_dmem_data_out [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[30]_i_1 
       (.I0(\processor/mem_rd_data [30]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [30]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [30]),
        .O(\processor/ex_dmem_data_out [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[31]_i_1 
       (.I0(\processor/mem_rd_data [31]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [31]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [31]),
        .O(\processor/ex_dmem_data_out [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0082000000000082)) 
    \dmem_data_out_p[31]_i_2 
       (.I0(\dmem_data_out_p[31]_i_4_n_0 ),
        .I1(\processor/execute/rs2_addr [4]),
        .I2(\processor/mem_rd_address [4]),
        .I3(\dmem_data_out_p[31]_i_5_n_0 ),
        .I4(\processor/mem_rd_address [3]),
        .I5(\processor/execute/rs2_addr [3]),
        .O(\dmem_data_out_p[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2002000000002002)) 
    \dmem_data_out_p[31]_i_3 
       (.I0(\dmem_data_out_p[31]_i_6_n_0 ),
        .I1(\dmem_data_out_p[31]_i_7_n_0 ),
        .I2(\processor/execute/rs2_addr [3]),
        .I3(\processor/wb_rd_address [3]),
        .I4(\processor/execute/rs2_addr [4]),
        .I5(\processor/wb_rd_address [4]),
        .O(\dmem_data_out_p[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAA8)) 
    \dmem_data_out_p[31]_i_4 
       (.I0(\processor/mem_rd_write ),
        .I1(\processor/mem_rd_address [2]),
        .I2(\processor/mem_rd_address [4]),
        .I3(\processor/mem_rd_address [1]),
        .I4(\processor/mem_rd_address [0]),
        .I5(\processor/mem_rd_address [3]),
        .O(\dmem_data_out_p[31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    \dmem_data_out_p[31]_i_5 
       (.I0(\processor/mem_rd_address [1]),
        .I1(\processor/execute/rs2_addr [1]),
        .I2(\processor/mem_rd_address [2]),
        .I3(\processor/execute/rs2_addr [2]),
        .I4(\processor/execute/rs2_addr [0]),
        .I5(\processor/mem_rd_address [0]),
        .O(\dmem_data_out_p[31]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAA8)) 
    \dmem_data_out_p[31]_i_6 
       (.I0(\processor/wb_rd_write ),
        .I1(\processor/wb_rd_address [2]),
        .I2(\processor/wb_rd_address [4]),
        .I3(\processor/wb_rd_address [1]),
        .I4(\processor/wb_rd_address [0]),
        .I5(\processor/wb_rd_address [3]),
        .O(\dmem_data_out_p[31]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    \dmem_data_out_p[31]_i_7 
       (.I0(\processor/execute/rs2_addr [2]),
        .I1(\processor/wb_rd_address [2]),
        .I2(\processor/wb_rd_address [1]),
        .I3(\processor/execute/rs2_addr [1]),
        .I4(\processor/wb_rd_address [0]),
        .I5(\processor/execute/rs2_addr [0]),
        .O(\dmem_data_out_p[31]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[3]_i_1 
       (.I0(\processor/mem_rd_data [3]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [3]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [3]),
        .O(\processor/ex_dmem_data_out [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[4]_i_1 
       (.I0(\processor/mem_rd_data [4]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [4]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [4]),
        .O(\processor/ex_dmem_data_out [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[5]_i_1 
       (.I0(\processor/mem_rd_data [5]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [5]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [5]),
        .O(\processor/ex_dmem_data_out [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[6]_i_1 
       (.I0(\processor/mem_rd_data [6]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [6]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [6]),
        .O(\processor/ex_dmem_data_out [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[7]_i_1 
       (.I0(\processor/mem_rd_data[7]_repN_1 ),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [7]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [7]),
        .O(\processor/ex_dmem_data_out [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[8]_i_1 
       (.I0(\processor/mem_rd_data [8]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [8]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [8]),
        .O(\processor/ex_dmem_data_out [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCAA00AAFFFFFFFF)) 
    \dmem_data_out_p[8]_i_2 
       (.I0(rd_data[8]),
        .I1(\mem_size[0]_repN ),
        .I2(\mem_size[1]_repN ),
        .I3(\rd_data_out[31]_i_4_n_0 ),
        .I4(\dmem_if/dmem_data_out_reg_n_0_[8] ),
        .I5(\rd_data_out[15]_i_3_n_0 ),
        .O(\processor/mem_rd_data [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dmem_data_out_p[9]_i_1 
       (.I0(\processor/mem_rd_data [9]),
        .I1(\dmem_data_out_p[31]_i_2_n_0 ),
        .I2(\processor/wb_rd_data [9]),
        .I3(\dmem_data_out_p[31]_i_3_n_0 ),
        .I4(\processor/rs2_data [9]),
        .O(\processor/ex_dmem_data_out [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCAA00AAFFFFFFFF)) 
    \dmem_data_out_p[9]_i_2 
       (.I0(rd_data[9]),
        .I1(\mem_size[0]_repN ),
        .I2(\mem_size[1]_repN ),
        .I3(\rd_data_out[31]_i_4_n_0 ),
        .I4(\dmem_if/dmem_data_out_reg_n_0_[9] ),
        .I5(\rd_data_out[15]_i_3_n_0 ),
        .O(\processor/mem_rd_data [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \dmem_data_size_p[0]_i_1 
       (.I0(\processor/ex_dmem_data_size [1]),
        .I1(\processor/ex_mem_size ),
        .O(\processor/ex_dmem_data_size [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000020000000)) 
    \dmem_if/dmem_data_out[31]_i_1 
       (.I0(\dmem_data_out[23]_i_3_n_0 ),
        .I1(reset),
        .I2(\dmem_if/state_reg_n_0_ ),
        .I3(\arbiter/state [1]),
        .I4(wb_ack_in),
        .I5(\arbiter/state [0]),
        .O(\dmem_if/dmem_data_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[0] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[0]),
        .Q(\dmem_if/dmem_data_out_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[10] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[10]),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[11] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[11]),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[12] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[12]),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[13] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[13]),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[14] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[14]),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[15] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[15]),
        .Q(p_1_in0),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[16] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[16]),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[17] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[17]),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[18] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[18]),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[19] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[19]),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[1] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[1]),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[20] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[20]),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[21] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[21]),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[22] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[22]),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[23] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[23]),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[24] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(\dmem_data_out[24]_i_1_n_0 ),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[24] ),
        .R(\dmem_if/dmem_data_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[25] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(\dmem_data_out[25]_i_1_n_0 ),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[25] ),
        .R(\dmem_if/dmem_data_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[26] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(\dmem_data_out[26]_i_1_n_0 ),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[26] ),
        .R(\dmem_if/dmem_data_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[27] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(\dmem_data_out[27]_i_1_n_0 ),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[27] ),
        .R(\dmem_if/dmem_data_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[28] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(\dmem_data_out[28]_i_1_n_0 ),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[28] ),
        .R(\dmem_if/dmem_data_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[29] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(\dmem_data_out[29]_i_1_n_0 ),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[29] ),
        .R(\dmem_if/dmem_data_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[2] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[2]),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[30] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(\dmem_data_out[30]_i_1_n_0 ),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[30] ),
        .R(\dmem_if/dmem_data_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[31] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(\dmem_data_out[31]_i_2_n_0 ),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[31] ),
        .R(\dmem_if/dmem_data_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[3] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[3]),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[4] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[4]),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[5] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[5]),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[6] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[6]),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[7] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[7]),
        .Q(p_0_in0),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "dmem_if/dmem_data_out_reg[7]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[7]_replica 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[7]),
        .Q(p_0_in0_repN),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[8] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[8]),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_data_out_reg[9] 
       (.C(clk),
        .CE(\dmem_data_out[23]_i_1_n_0 ),
        .D(SHIFT_RIGHT[9]),
        .Q(\dmem_if/dmem_data_out_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/dmem_r_ack_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(dmem_r_ack_i_1_n_0),
        .Q(dmem_read_ack),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair65" *) 
  LUT4 #(
    .INIT(16'h0F10)) 
    \dmem_if/state[0]_i_1 
       (.I0(dmem_write_req),
        .I1(\dmem_if/state_reg_n_0_[1] ),
        .I2(\state[1]_i_3_n_0 ),
        .I3(\dmem_if/state_reg_n_0_ ),
        .O(\dmem_if/state ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair65" *) 
  LUT4 #(
    .INIT(16'h0F20)) 
    \dmem_if/state[1]_i_1 
       (.I0(dmem_write_req),
        .I1(\dmem_if/state_reg_n_0_ ),
        .I2(\state[1]_i_3_n_0 ),
        .I3(\dmem_if/state_reg_n_0_[1] ),
        .O(\dmem_if/state[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/state_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\dmem_if/state ),
        .Q(\dmem_if/state_reg_n_0_ ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/state_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\dmem_if/state[1]_i_1_n_0 ),
        .Q(\dmem_if/state_reg_n_0_[1] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][0] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address[0]),
        .Q(\dmem_if_outputs[adr] [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][10] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[10]),
        .Q(\dmem_if_outputs[adr] [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][11] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[11]),
        .Q(\dmem_if_outputs[adr] [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][12] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[12]),
        .Q(\dmem_if_outputs[adr] [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][13] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[13]),
        .Q(\dmem_if_outputs[adr] [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][14] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[14]),
        .Q(\dmem_if_outputs[adr] [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][15] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[15]),
        .Q(\dmem_if_outputs[adr] [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][16] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[16]),
        .Q(\dmem_if_outputs[adr] [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][17] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[17]),
        .Q(\dmem_if_outputs[adr] [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][18] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[18]),
        .Q(\dmem_if_outputs[adr] [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][19] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[19]),
        .Q(\dmem_if_outputs[adr] [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][1] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address[1]),
        .Q(\dmem_if_outputs[adr] [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][20] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[20]),
        .Q(\dmem_if_outputs[adr] [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][21] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[21]),
        .Q(\dmem_if_outputs[adr] [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][22] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[22]),
        .Q(\dmem_if_outputs[adr] [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][23] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[23]),
        .Q(\dmem_if_outputs[adr] [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][24] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[24]),
        .Q(\dmem_if_outputs[adr] [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][25] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[25]),
        .Q(\dmem_if_outputs[adr] [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][26] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[26]),
        .Q(\dmem_if_outputs[adr] [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][27] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[27]),
        .Q(\dmem_if_outputs[adr] [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][28] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[28]),
        .Q(\dmem_if_outputs[adr] [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][29] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[29]),
        .Q(\dmem_if_outputs[adr] [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][2] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[2]),
        .Q(\dmem_if_outputs[adr] [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][30] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[30]),
        .Q(\dmem_if_outputs[adr] [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][31] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[31]),
        .Q(\dmem_if_outputs[adr] [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][3] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[3]),
        .Q(\dmem_if_outputs[adr] [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][4] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[4]),
        .Q(\dmem_if_outputs[adr] [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][5] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[5]),
        .Q(\dmem_if_outputs[adr] [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][6] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[6]),
        .Q(\dmem_if_outputs[adr] [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][7] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[7]),
        .Q(\dmem_if_outputs[adr] [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][8] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[8]),
        .Q(\dmem_if_outputs[adr] [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[adr][9] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(dmem_address__0[9]),
        .Q(\dmem_if_outputs[adr] [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[cyc] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\wb_outputs[cyc]_i_1_n_0 ),
        .Q(dmem_if_outputs),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][0] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(\wb_outputs[dat][0]_i_1_n_0 ),
        .Q(\dmem_if_outputs[dat] [0]),
        .R(\wb_outputs[dat][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][10] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(SHIFT_LEFT[10]),
        .Q(\dmem_if_outputs[dat] [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][11] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(SHIFT_LEFT[11]),
        .Q(\dmem_if_outputs[dat] [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][12] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(SHIFT_LEFT[12]),
        .Q(\dmem_if_outputs[dat] [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][13] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(SHIFT_LEFT[13]),
        .Q(\dmem_if_outputs[dat] [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][14] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(SHIFT_LEFT[14]),
        .Q(\dmem_if_outputs[dat] [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][15] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(SHIFT_LEFT[15]),
        .Q(\dmem_if_outputs[dat] [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][16] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(SHIFT_LEFT[16]),
        .Q(\dmem_if_outputs[dat] [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][17] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(SHIFT_LEFT[17]),
        .Q(\dmem_if_outputs[dat] [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][18] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(SHIFT_LEFT[18]),
        .Q(\dmem_if_outputs[dat] [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][19] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(SHIFT_LEFT[19]),
        .Q(\dmem_if_outputs[dat] [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][1] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(\wb_outputs[dat][1]_i_1_n_0 ),
        .Q(\dmem_if_outputs[dat] [1]),
        .R(\wb_outputs[dat][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][20] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(SHIFT_LEFT[20]),
        .Q(\dmem_if_outputs[dat] [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][21] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(SHIFT_LEFT[21]),
        .Q(\dmem_if_outputs[dat] [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][22] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(SHIFT_LEFT[22]),
        .Q(\dmem_if_outputs[dat] [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][23] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(SHIFT_LEFT[23]),
        .Q(\dmem_if_outputs[dat] [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][24] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(SHIFT_LEFT[24]),
        .Q(\dmem_if_outputs[dat] [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][25] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(SHIFT_LEFT[25]),
        .Q(\dmem_if_outputs[dat] [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][26] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(SHIFT_LEFT[26]),
        .Q(\dmem_if_outputs[dat] [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][27] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(SHIFT_LEFT[27]),
        .Q(\dmem_if_outputs[dat] [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][28] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(SHIFT_LEFT[28]),
        .Q(\dmem_if_outputs[dat] [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][29] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(SHIFT_LEFT[29]),
        .Q(\dmem_if_outputs[dat] [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][2] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(\wb_outputs[dat][2]_i_1_n_0 ),
        .Q(\dmem_if_outputs[dat] [2]),
        .R(\wb_outputs[dat][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][30] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(SHIFT_LEFT[30]),
        .Q(\dmem_if_outputs[dat] [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][31] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(SHIFT_LEFT[31]),
        .Q(\dmem_if_outputs[dat] [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][3] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(\wb_outputs[dat][3]_i_1_n_0 ),
        .Q(\dmem_if_outputs[dat] [3]),
        .R(\wb_outputs[dat][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][4] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(\wb_outputs[dat][4]_i_1_n_0 ),
        .Q(\dmem_if_outputs[dat] [4]),
        .R(\wb_outputs[dat][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][5] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(\wb_outputs[dat][5]_i_1_n_0 ),
        .Q(\dmem_if_outputs[dat] [5]),
        .R(\wb_outputs[dat][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][6] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(\wb_outputs[dat][6]_i_1_n_0 ),
        .Q(\dmem_if_outputs[dat] [6]),
        .R(\wb_outputs[dat][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][7] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(\wb_outputs[dat][7]_i_2_n_0 ),
        .Q(\dmem_if_outputs[dat] [7]),
        .R(\wb_outputs[dat][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][8] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(SHIFT_LEFT[8]),
        .Q(\dmem_if_outputs[dat] [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[dat][9] 
       (.C(clk),
        .CE(\wb_outputs[dat][31]_i_1_n_0 ),
        .D(SHIFT_LEFT[9]),
        .Q(\dmem_if_outputs[dat] [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[sel][0] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(\wb_outputs[sel][0]_i_1_n_0 ),
        .Q(\dmem_if_outputs[sel] [0]),
        .S(\wb_outputs[sel][3]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[sel][1] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(\wb_outputs[sel][1]_i_1_n_0 ),
        .Q(\dmem_if_outputs[sel] [1]),
        .S(\wb_outputs[sel][3]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[sel][2] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(\wb_outputs[sel][2]_i_1_n_0 ),
        .Q(\dmem_if_outputs[sel] [2]),
        .S(\wb_outputs[sel][3]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[sel][3] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1_n_0 ),
        .D(\wb_outputs[sel][3]_i_2_n_0 ),
        .Q(\dmem_if_outputs[sel] [3]),
        .S(\wb_outputs[sel][3]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \dmem_if/wb_outputs_reg[we] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\wb_outputs[we]_i_1_n_0 ),
        .Q(\dmem_if_outputs[we] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFAAAA10000000)) 
    dmem_r_ack_i_1
       (.I0(\dmem_if/state_reg_n_0_[1] ),
        .I1(\arbiter/state [0]),
        .I2(wb_ack_in),
        .I3(\arbiter/state [1]),
        .I4(\dmem_if/state_reg_n_0_ ),
        .I5(dmem_read_ack),
        .O(dmem_r_ack_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    dmem_read_req_p_i_1
       (.I0(\processor/ex_mem_op [2]),
        .I1(\processor/ex_mem_op [1]),
        .I2(\mem_op[2]_i_5_n_0 ),
        .O(\processor/ex_dmem_read_req ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    dmem_write_req_p_i_1
       (.I0(\processor/ex_mem_op [0]),
        .I1(\processor/ex_mem_op [2]),
        .I2(\processor/ex_mem_op [1]),
        .I3(\mem_op[2]_i_5_n_0 ),
        .O(\processor/ex_dmem_write_req ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0FFF00F008FB08FB)) 
    \exception_context_out[badaddr][0]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [0]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\mem_op[2]_i_5_n_0 ),
        .I3(exception_context_out),
        .I4(\processor/mem_exception_context[badaddr] [0]),
        .I5(\processor/mem_exception ),
        .O(\processor/ex_exception_context[badaddr] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00D700FF)) 
    \exception_context_out[badaddr][0]_i_2 
       (.I0(\processor/ex_rd_data [0]),
        .I1(\processor/ex_dmem_data_size [1]),
        .I2(\processor/ex_mem_size ),
        .I3(\exception_context_out[badaddr][1]_i_4_n_0 ),
        .I4(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .O(exception_context_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][10]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [10]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [10]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][10]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][10]_i_2 
       (.I0(\processor/ex_rd_data [10]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[10]_i_2_n_0 ),
        .O(\exception_context_out[badaddr][10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][11]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [11]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [11]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][11]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][11]_i_2 
       (.I0(\processor/ex_rd_data [11]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[11]_i_2_n_0 ),
        .O(\exception_context_out[badaddr][11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][12]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [12]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [12]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][12]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][12]_i_2 
       (.I0(\processor/ex_rd_data [12]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[12]_i_3_n_0 ),
        .O(\exception_context_out[badaddr][12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][13]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [13]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [13]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][13]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][13]_i_2 
       (.I0(\processor/ex_rd_data [13]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[13]_i_2_n_0 ),
        .O(\exception_context_out[badaddr][13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][14]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [14]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [14]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][14]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][14]_i_2 
       (.I0(\processor/ex_rd_data [14]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[14]_i_2_n_0 ),
        .O(\exception_context_out[badaddr][14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][15]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [15]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [15]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][15]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][15]_i_2 
       (.I0(\processor/ex_rd_data [15]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[15]_i_2_n_0 ),
        .O(\exception_context_out[badaddr][15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][16]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [16]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [16]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][16]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][16]_i_2 
       (.I0(\processor/ex_rd_data [16]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[16]_i_3_n_0 ),
        .O(\exception_context_out[badaddr][16]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][17]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [17]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [17]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][17]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][17]_i_2 
       (.I0(\processor/ex_rd_data [17]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[17]_i_2_n_0 ),
        .O(\exception_context_out[badaddr][17]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][18]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [18]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [18]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][18]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][18]_i_2 
       (.I0(\processor/ex_rd_data [18]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[18]_i_2_n_0 ),
        .O(\exception_context_out[badaddr][18]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][19]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [19]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [19]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][19]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][19]_i_2 
       (.I0(\processor/ex_rd_data [19]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[19]_i_2_n_0 ),
        .O(\exception_context_out[badaddr][19]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0FFF00F008FB08FB)) 
    \exception_context_out[badaddr][1]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [1]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\mem_op[2]_i_5_n_0 ),
        .I3(\exception_context_out[badaddr][1]_i_2_n_0 ),
        .I4(\processor/mem_exception_context[badaddr] [1]),
        .I5(\processor/mem_exception ),
        .O(\processor/ex_exception_context[badaddr] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAA0A2AAA)) 
    \exception_context_out[badaddr][1]_i_2 
       (.I0(\exception_context_out[badaddr][1]_i_3_n_0_repN ),
        .I1(\processor/ex_rd_data [0]),
        .I2(\processor/ex_rd_data [1]),
        .I3(\processor/ex_dmem_data_size [1]),
        .I4(\processor/ex_mem_size ),
        .I5(\exception_context_out[badaddr][1]_i_4_n_0 ),
        .O(\exception_context_out[badaddr][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "exception_context_out[badaddr][1]_i_3" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \exception_context_out[badaddr][1]_i_3_replica 
       (.I0(\pc[1]_i_3_n_0 ),
        .I1(\mem_op[2]_i_4_n_0 ),
        .O(\exception_context_out[badaddr][1]_i_3_n_0_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h2)) 
    \exception_context_out[badaddr][1]_i_3_rewire 
       (.I0(\pc[1]_i_3_n_0 ),
        .O(\exception_context_out[badaddr][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \exception_context_out[badaddr][1]_i_4 
       (.I0(\mem_op[2]_i_4_n_0 ),
        .I1(\pc[0]_i_3_n_0 ),
        .O(\exception_context_out[badaddr][1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][20]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [20]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [20]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][20]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][20]_i_2 
       (.I0(\processor/ex_rd_data [20]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[20]_i_3_n_0 ),
        .O(\exception_context_out[badaddr][20]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][21]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [21]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [21]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][21]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][21]_i_2 
       (.I0(\processor/ex_rd_data [21]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[21]_i_2_n_0 ),
        .O(\exception_context_out[badaddr][21]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][22]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [22]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [22]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][22]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][22]_i_2 
       (.I0(\processor/ex_rd_data [22]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[22]_i_2_n_0 ),
        .O(\exception_context_out[badaddr][22]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][23]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [23]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [23]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][23]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][23]_i_2 
       (.I0(\processor/ex_rd_data [23]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[23]_i_2_n_0 ),
        .O(\exception_context_out[badaddr][23]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][24]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [24]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [24]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][24]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][24]_i_2 
       (.I0(\processor/ex_rd_data [24]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[24]_i_3_n_0 ),
        .O(\exception_context_out[badaddr][24]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][25]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [25]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [25]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][25]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][25]_i_2 
       (.I0(\processor/ex_rd_data [25]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[25]_i_2_n_0 ),
        .O(\exception_context_out[badaddr][25]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][26]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [26]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [26]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][26]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][26]_i_2 
       (.I0(\processor/ex_rd_data [26]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[26]_i_2_n_0 ),
        .O(\exception_context_out[badaddr][26]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][27]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [27]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [27]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][27]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][27]_i_2 
       (.I0(\processor/ex_rd_data [27]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[27]_i_2_n_0 ),
        .O(\exception_context_out[badaddr][27]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][28]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [28]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [28]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][28]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][28]_i_2 
       (.I0(\processor/ex_rd_data [28]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[28]_i_3_n_0 ),
        .O(\exception_context_out[badaddr][28]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][29]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [29]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [29]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][29]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][29]_i_2 
       (.I0(\processor/ex_rd_data [29]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[29]_i_2_n_0 ),
        .O(\exception_context_out[badaddr][29]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][2]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [2]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [2]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][2]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][2]_i_2 
       (.I0(\processor/ex_rd_data [2]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[2]_i_3_n_0 ),
        .O(\exception_context_out[badaddr][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][30]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [30]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [30]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][30]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][30]_i_2 
       (.I0(\processor/ex_rd_data [30]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[30]_i_2_n_0 ),
        .O(\exception_context_out[badaddr][30]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \exception_context_out[badaddr][31]_i_1 
       (.I0(\mem_op[2]_i_5_n_0 ),
        .I1(reset),
        .O(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][31]_i_2 
       (.I0(\processor/wb_exception_context[badaddr] [31]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [31]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][31]_i_4_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \exception_context_out[badaddr][31]_i_3 
       (.I0(\processor/wb_exception ),
        .I1(\exception_context_out[ie1]_i_4_n_0 ),
        .O(\exception_context_out[badaddr][31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][31]_i_4 
       (.I0(\processor/ex_rd_data [31]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[31]_i_4_n_0 ),
        .O(\exception_context_out[badaddr][31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hC7D7)) 
    \exception_context_out[badaddr][31]_i_5 
       (.I0(\processor/ex_rd_data [0]),
        .I1(\processor/ex_dmem_data_size [1]),
        .I2(\processor/ex_mem_size ),
        .I3(\processor/ex_rd_data [1]),
        .O(\exception_context_out[badaddr][31]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h0D)) 
    \exception_context_out[badaddr][31]_i_6_rewire 
       (.I0(\mem_op[2]_i_4_n_0 ),
        .I1(\exception_context_out[badaddr][1]_i_3_n_0 ),
        .I2(\exception_context_out[badaddr][1]_i_4_n_0 ),
        .O(\exception_context_out[badaddr][31]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][3]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [3]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [3]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][3]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][3]_i_2 
       (.I0(\processor/ex_rd_data [3]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[3]_i_3_n_0 ),
        .O(\exception_context_out[badaddr][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][4]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [4]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [4]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][4]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][4]_i_2 
       (.I0(\processor/ex_rd_data [4]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[4]_i_2_n_0 ),
        .O(\exception_context_out[badaddr][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][5]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [5]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [5]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][5]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][5]_i_2 
       (.I0(\processor/ex_rd_data [5]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[5]_i_2_n_0 ),
        .O(\exception_context_out[badaddr][5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][6]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [6]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [6]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][6]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][6]_i_2 
       (.I0(\processor/ex_rd_data [6]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[6]_i_2_n_0 ),
        .O(\exception_context_out[badaddr][6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][7]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [7]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [7]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][7]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][7]_i_2 
       (.I0(\processor/ex_rd_data [7]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[7]_i_2_n_0 ),
        .O(\exception_context_out[badaddr][7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][8]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [8]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [8]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][8]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][8]_i_2 
       (.I0(\processor/ex_rd_data [8]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[8]_i_2_n_0 ),
        .O(\exception_context_out[badaddr][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[badaddr][9]_i_1 
       (.I0(\processor/wb_exception_context[badaddr] [9]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [9]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[badaddr][9]_i_2_n_0 ),
        .O(\processor/ex_exception_context[badaddr] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \exception_context_out[badaddr][9]_i_2 
       (.I0(\processor/ex_rd_data [9]),
        .I1(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I3(\pc[9]_i_2_n_0 ),
        .O(\exception_context_out[badaddr][9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00FF00AAAACFC0)) 
    \exception_context_out[cause][0]_i_1 
       (.I0(\processor/mem_exception_context[cause] [0]),
        .I1(\processor/wb_exception_context[cause] [0]),
        .I2(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I3(\exception_context_out[cause][0]_i_2_n_0 ),
        .I4(\processor/mem_exception ),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\processor/ex_exception_context[cause] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \exception_context_out[cause][0]_i_10 
       (.I0(irq[7]),
        .I1(\processor/execute/mie [31]),
        .I2(\exception_context_out[cause][0]_i_7_n_0 ),
        .I3(\processor/wb_csr_data [31]),
        .I4(\exception_context_out[cause][0]_i_8_n_0 ),
        .I5(\processor/mem_csr_data [31]),
        .O(\exception_context_out[cause][0]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAA8A8000008A80)) 
    \exception_context_out[cause][0]_i_11 
       (.I0(irq[5]),
        .I1(\processor/wb_csr_data [29]),
        .I2(\exception_context_out[cause][0]_i_7_n_0 ),
        .I3(\processor/execute/mie [29]),
        .I4(\exception_context_out[cause][0]_i_8_n_0 ),
        .I5(\processor/mem_csr_data [29]),
        .O(\exception_context_out[cause][0]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \exception_context_out[cause][0]_i_12 
       (.I0(irq[4]),
        .I1(\processor/execute/mie [28]),
        .I2(\exception_context_out[cause][0]_i_7_n_0 ),
        .I3(\processor/wb_csr_data [28]),
        .I4(\exception_context_out[cause][0]_i_8_n_0 ),
        .I5(\processor/mem_csr_data [28]),
        .O(\exception_context_out[cause][0]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \exception_context_out[cause][0]_i_13 
       (.I0(irq[3]),
        .I1(\processor/execute/mie [27]),
        .I2(\exception_context_out[cause][0]_i_7_n_0 ),
        .I3(\processor/wb_csr_data [27]),
        .I4(\exception_context_out[cause][0]_i_8_n_0 ),
        .I5(\processor/mem_csr_data [27]),
        .O(\exception_context_out[cause][0]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \exception_context_out[cause][0]_i_14 
       (.I0(irq[2]),
        .I1(\processor/execute/mie [26]),
        .I2(\exception_context_out[cause][0]_i_7_n_0 ),
        .I3(\processor/wb_csr_data [26]),
        .I4(\exception_context_out[cause][0]_i_8_n_0 ),
        .I5(\processor/mem_csr_data [26]),
        .O(\exception_context_out[cause][0]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \exception_context_out[cause][0]_i_15 
       (.I0(\processor/mem_csr_address [1]),
        .I1(\processor/mem_csr_address [7]),
        .O(\exception_context_out[cause][0]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0E000000)) 
    \exception_context_out[cause][0]_i_16 
       (.I0(\processor/mem_csr_write [0]),
        .I1(\processor/mem_csr_write [1]),
        .I2(\processor/mem_csr_address[4]_repN_1 ),
        .I3(\processor/mem_csr_address [8]),
        .I4(\processor/mem_csr_address [2]),
        .O(\exception_context_out[cause][0]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \exception_context_out[cause][0]_i_17 
       (.I0(\processor/mem_csr_address [11]),
        .I1(\processor/mem_csr_address [3]),
        .I2(\processor/mem_csr_address [10]),
        .I3(\processor/mem_csr_address [0]),
        .O(\exception_context_out[cause][0]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h54545454000000FF)) 
    \exception_context_out[cause][0]_i_2 
       (.I0(\exception_context_out[cause][0]_i_3_n_0 ),
        .I1(\exception_context_out[cause][0]_i_4_n_0 ),
        .I2(\exception_context_out[cause][0]_i_5_n_0 ),
        .I3(\exception_context_out[cause][0]_i_6_n_0 ),
        .I4(\exception_context_out[cause][5]_i_3_n_0 ),
        .I5(\exception_context_out[cause][5]_i_4_n_0 ),
        .O(\exception_context_out[cause][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAA8A8000008A80)) 
    \exception_context_out[cause][0]_i_3 
       (.I0(irq[0]),
        .I1(\processor/wb_csr_data [24]),
        .I2(\exception_context_out[cause][0]_i_7_n_0 ),
        .I3(\processor/execute/mie [24]),
        .I4(\exception_context_out[cause][0]_i_8_n_0 ),
        .I5(\processor/mem_csr_data [24]),
        .O(\exception_context_out[cause][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAA8A8000008A80)) 
    \exception_context_out[cause][0]_i_4 
       (.I0(irq[1]),
        .I1(\processor/wb_csr_data [25]),
        .I2(\exception_context_out[cause][0]_i_7_n_0 ),
        .I3(\processor/execute/mie [25]),
        .I4(\exception_context_out[cause][0]_i_8_n_0 ),
        .I5(\processor/mem_csr_data [25]),
        .O(\exception_context_out[cause][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFF00F1)) 
    \exception_context_out[cause][0]_i_5 
       (.I0(\exception_context_out[cause][0]_i_9_n_0 ),
        .I1(\exception_context_out[cause][0]_i_10_n_0 ),
        .I2(\exception_context_out[cause][0]_i_11_n_0 ),
        .I3(\exception_context_out[cause][0]_i_12_n_0 ),
        .I4(\exception_context_out[cause][0]_i_13_n_0 ),
        .I5(\exception_context_out[cause][0]_i_14_n_0 ),
        .O(\exception_context_out[cause][0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h002A)) 
    \exception_context_out[cause][0]_i_6 
       (.I0(\exception_context_out[cause][4]_i_3_n_0 ),
        .I1(\processor/execute/decode_exception ),
        .I2(\processor/execute/decode_exception_cause [0]),
        .I3(\exception_context_out[cause][5]_i_5_n_0 ),
        .O(\exception_context_out[cause][0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \exception_context_out[cause][0]_i_7 
       (.I0(\exception_context_out[ie1]_i_10_n_0 ),
        .I1(\processor/wb_csr_address [2]),
        .I2(\exception_context_out[ie1]_i_11_n_0 ),
        .O(\exception_context_out[cause][0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000001000000)) 
    \exception_context_out[cause][0]_i_8 
       (.I0(\processor/mem_csr_address [6]),
        .I1(\processor/mem_csr_address [5]),
        .I2(\exception_context_out[cause][0]_i_15_n_0 ),
        .I3(\exception_context_out[cause][0]_i_16_n_0 ),
        .I4(\processor/mem_csr_address [9]),
        .I5(\exception_context_out[cause][0]_i_17_n_0 ),
        .O(\exception_context_out[cause][0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \exception_context_out[cause][0]_i_9 
       (.I0(irq[6]),
        .I1(\processor/execute/mie [30]),
        .I2(\exception_context_out[cause][0]_i_7_n_0 ),
        .I3(\processor/wb_csr_data [30]),
        .I4(\exception_context_out[cause][0]_i_8_n_0 ),
        .I5(\processor/mem_csr_data [30]),
        .O(\exception_context_out[cause][0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000F088FFFFF0BB)) 
    \exception_context_out[cause][1]_i_1 
       (.I0(\processor/wb_exception_context[cause] [1]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[cause] [1]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[cause][1]_i_2_n_0 ),
        .O(\processor/ex_exception_context[cause] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFF08AA)) 
    \exception_context_out[cause][1]_i_2 
       (.I0(\exception_context_out[cause][1]_i_3_n_0 ),
        .I1(\exception_context_out[cause][3]_i_4_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I3(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I4(\exception_context_out[cause][5]_i_2_n_0 ),
        .I5(\exception_context_out[cause][1]_i_4_n_0 ),
        .O(\exception_context_out[cause][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5455)) 
    \exception_context_out[cause][1]_i_3 
       (.I0(\processor/execute/decode_exception ),
        .I1(\processor/ex_mem_op [2]),
        .I2(\processor/ex_mem_op [1]),
        .I3(\processor/ex_mem_op [0]),
        .O(\exception_context_out[cause][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0010101000100010)) 
    \exception_context_out[cause][1]_i_4 
       (.I0(\exception_context_out[cause][0]_i_3_n_0 ),
        .I1(\exception_context_out[cause][0]_i_4_n_0 ),
        .I2(\processor/ex_exception_context[ie] ),
        .I3(\exception_context_out[cause][2]_i_8_n_0 ),
        .I4(\exception_context_out[cause][2]_i_7_n_0 ),
        .I5(\exception_context_out[cause][2]_i_6_n_0 ),
        .O(\exception_context_out[cause][1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000F088FFFFF0BB)) 
    \exception_context_out[cause][2]_i_1 
       (.I0(\processor/wb_exception_context[cause] [2]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[cause] [2]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[cause][2]_i_2_n_0 ),
        .O(\processor/ex_exception_context[cause] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF2F2F2F2F200F2F2)) 
    \exception_context_out[cause][2]_i_2 
       (.I0(\exception_context_out[cause][3]_i_6_n_0 ),
        .I1(\exception_context_out[cause][2]_i_3_n_0 ),
        .I2(\exception_context_out[cause][5]_i_2_n_0 ),
        .I3(\exception_context_out[cause][2]_i_4_n_0 ),
        .I4(\processor/ex_exception_context[ie] ),
        .I5(\exception_context_out[cause][2]_i_5_n_0 ),
        .O(\exception_context_out[cause][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \exception_context_out[cause][2]_i_3 
       (.I0(\processor/execute/decode_exception ),
        .I1(\processor/execute/decode_exception_cause [2]),
        .O(\exception_context_out[cause][2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \exception_context_out[cause][2]_i_4 
       (.I0(\exception_context_out[cause][2]_i_6_n_0 ),
        .I1(\exception_context_out[cause][2]_i_7_n_0 ),
        .O(\exception_context_out[cause][2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEF)) 
    \exception_context_out[cause][2]_i_5 
       (.I0(\exception_context_out[cause][0]_i_3_n_0 ),
        .I1(\exception_context_out[cause][0]_i_4_n_0 ),
        .I2(\exception_context_out[cause][2]_i_8_n_0 ),
        .O(\exception_context_out[cause][2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \exception_context_out[cause][2]_i_6 
       (.I0(\exception_context_out[cause][0]_i_9_n_0 ),
        .I1(\exception_context_out[cause][0]_i_10_n_0 ),
        .O(\exception_context_out[cause][2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \exception_context_out[cause][2]_i_7 
       (.I0(\exception_context_out[cause][0]_i_12_n_0 ),
        .I1(\exception_context_out[cause][0]_i_11_n_0 ),
        .O(\exception_context_out[cause][2]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \exception_context_out[cause][2]_i_8 
       (.I0(\exception_context_out[cause][0]_i_14_n_0 ),
        .I1(\exception_context_out[cause][0]_i_13_n_0 ),
        .O(\exception_context_out[cause][2]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00C5FFC500C500C5)) 
    \exception_context_out[cause][3]_i_1 
       (.I0(\exception_context_out[cause][3]_i_2_n_0 ),
        .I1(\processor/mem_exception_context[cause] [3]),
        .I2(\processor/mem_exception ),
        .I3(\mem_op[2]_i_5_n_0 ),
        .I4(\exception_context_out[cause][5]_i_2_n_0 ),
        .I5(\exception_context_out[cause][3]_i_3_n_0 ),
        .O(\processor/ex_exception_context[cause] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5C5F5F5F5C5C5C5C)) 
    \exception_context_out[cause][3]_i_2 
       (.I0(\processor/wb_exception_context[cause] [3]),
        .I1(\exception_context_out[cause][5]_i_2_n_0 ),
        .I2(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I3(\processor/execute/decode_exception_cause [3]),
        .I4(\processor/execute/decode_exception ),
        .I5(\exception_context_out[cause][4]_i_3_n_0 ),
        .O(\exception_context_out[cause][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88888888FF88FF8F)) 
    \exception_context_out[cause][3]_i_3 
       (.I0(\processor/execute/decode_exception_cause [3]),
        .I1(\processor/execute/decode_exception ),
        .I2(\exception_context_out[cause][3]_i_4_n_0 ),
        .I3(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .I4(\exception_context_out[cause][3]_i_5_n_0 ),
        .I5(\exception_context_out[cause][3]_i_6_n_0 ),
        .O(\exception_context_out[cause][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \exception_context_out[cause][3]_i_4 
       (.I0(\processor/ex_mem_op [1]),
        .I1(\processor/ex_mem_op [2]),
        .O(\exception_context_out[cause][3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \exception_context_out[cause][3]_i_5 
       (.I0(\processor/ex_mem_op [1]),
        .I1(\processor/ex_mem_op [2]),
        .I2(\processor/ex_mem_op [0]),
        .O(\exception_context_out[cause][3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF555D)) 
    \exception_context_out[cause][3]_i_6 
       (.I0(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I1(\processor/ex_mem_op [0]),
        .I2(\processor/ex_mem_op [1]),
        .I3(\processor/ex_mem_op [2]),
        .I4(\processor/execute/decode_exception ),
        .O(\exception_context_out[cause][3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[cause][4]_i_1 
       (.I0(\processor/wb_exception_context[cause] [4]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[cause] [4]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[cause][4]_i_2_n_0 ),
        .O(\processor/ex_exception_context[cause] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAFBBB)) 
    \exception_context_out[cause][4]_i_2 
       (.I0(\exception_context_out[cause][5]_i_4_n_0 ),
        .I1(\exception_context_out[cause][4]_i_3_n_0 ),
        .I2(\processor/execute/decode_exception_cause [2]),
        .I3(\processor/execute/decode_exception ),
        .I4(\exception_context_out[cause][5]_i_5_n_0 ),
        .I5(\exception_context_out[cause][5]_i_3_n_0 ),
        .O(\exception_context_out[cause][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBBBBFBBBFFBFFB)) 
    \exception_context_out[cause][4]_i_3 
       (.I0(\processor/execute/decode_exception ),
        .I1(\exception_context_out[badaddr][31]_i_6_n_0 ),
        .I2(\processor/ex_mem_op [0]),
        .I3(\processor/ex_mem_op [2]),
        .I4(\processor/ex_mem_op [1]),
        .I5(\exception_context_out[badaddr][31]_i_5_n_0 ),
        .O(\exception_context_out[cause][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0BB0000F088)) 
    \exception_context_out[cause][5]_i_1 
       (.I0(\processor/wb_exception_context[cause] [5]),
        .I1(\exception_context_out[badaddr][31]_i_3_n_0 ),
        .I2(\processor/mem_exception_context[cause] [5]),
        .I3(\processor/mem_exception ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .I5(\exception_context_out[cause][5]_i_2_n_0 ),
        .O(\processor/ex_exception_context[cause] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \exception_context_out[cause][5]_i_2 
       (.I0(\exception_context_out[cause][5]_i_3_n_0 ),
        .I1(\exception_context_out[cause][5]_i_4_n_0 ),
        .I2(\exception_context_out[cause][5]_i_5_n_0 ),
        .O(\exception_context_out[cause][5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \exception_context_out[cause][5]_i_3 
       (.I0(\processor/ex_exception_context[ie] ),
        .I1(\exception_context_out[cause][5]_i_6_n_0 ),
        .O(\exception_context_out[cause][5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h8A)) 
    \exception_context_out[cause][5]_i_4 
       (.I0(\processor/ex_exception_context[ie] ),
        .I1(\exception_context_out[cause][2]_i_5_n_0 ),
        .I2(\exception_context_out[cause][2]_i_4_n_0 ),
        .O(\exception_context_out[cause][5]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \exception_context_out[cause][5]_i_5 
       (.I0(\processor/ex_exception_context[ie] ),
        .I1(\exception_context_out[cause][5]_i_7_n_0 ),
        .O(\exception_context_out[cause][5]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5555757FFFFF757F)) 
    \exception_context_out[cause][5]_i_6 
       (.I0(\processor/software_interrupt ),
        .I1(\processor/wb_csr_data [3]),
        .I2(\exception_context_out[cause][0]_i_7_n_0 ),
        .I3(\processor/execute/mie [3]),
        .I4(\exception_context_out[cause][5]_i_8_n_0 ),
        .I5(\processor/mem_csr_data [3]),
        .O(\exception_context_out[cause][5]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FF1D1DFFFFFFFF)) 
    \exception_context_out[cause][5]_i_7 
       (.I0(\processor/execute/mie [7]),
        .I1(\exception_context_out[cause][0]_i_7_n_0 ),
        .I2(\processor/wb_csr_data [7]),
        .I3(\processor/mem_csr_data [7]),
        .I4(\exception_context_out[cause][5]_i_8_n_0 ),
        .I5(\processor/timer_interrupt ),
        .O(\exception_context_out[cause][5]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002220)) 
    \exception_context_out[cause][5]_i_8 
       (.I0(\exception_context_out[cause][5]_i_9_n_0 ),
        .I1(\processor/mem_csr_address [4]),
        .I2(\processor/mem_csr_write [1]),
        .I3(\processor/mem_csr_write [0]),
        .I4(\exception_context_out[cause][0]_i_17_n_0 ),
        .O(\exception_context_out[cause][5]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000080000)) 
    \exception_context_out[cause][5]_i_9 
       (.I0(\processor/mem_csr_address [2]),
        .I1(\processor/mem_csr_address [9]),
        .I2(\processor/mem_csr_address [5]),
        .I3(\processor/mem_csr_address [6]),
        .I4(\processor/mem_csr_address [8]),
        .I5(\exception_context_out[cause][0]_i_15_n_0 ),
        .O(\exception_context_out[cause][5]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBABBBB888A8888)) 
    \exception_context_out[ie1]_i_1 
       (.I0(\processor/ex_exception_context[ie] ),
        .I1(\mem_op[2]_i_5_n_0 ),
        .I2(\processor/ex_branch [1]),
        .I3(\processor/ex_branch [0]),
        .I4(\processor/ex_branch [2]),
        .I5(\processor/ex_exception_context ),
        .O(\exception_context_out[ie1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \exception_context_out[ie1]_i_10 
       (.I0(\processor/wb_csr_address [8]),
        .I1(\processor/wb_csr_address [9]),
        .I2(\processor/wb_csr_address [10]),
        .I3(\processor/wb_csr_address [3]),
        .I4(\processor/wb_csr_address [11]),
        .I5(\processor/wb_csr_address [0]),
        .O(\exception_context_out[ie1]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFFFF)) 
    \exception_context_out[ie1]_i_11 
       (.I0(\processor/wb_csr_address [1]),
        .I1(\processor/wb_csr_address [7]),
        .I2(\processor/wb_csr_address [5]),
        .I3(\processor/wb_csr_address [6]),
        .I4(\processor/csr_unit/tohost_data1__0 ),
        .I5(\processor/wb_csr_address [4]),
        .O(\exception_context_out[ie1]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFE54BA10)) 
    \exception_context_out[ie1]_i_2 
       (.I0(\processor/mem_exception ),
        .I1(\exception_context_out[ie1]_i_4_n_0 ),
        .I2(\exception_context_out[ie1]_i_5_n_0 ),
        .I3(\processor/mem_exception_context[ie] ),
        .I4(\processor/mem_csr_data [0]),
        .O(\processor/ex_exception_context[ie] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFE54BA10)) 
    \exception_context_out[ie1]_i_3 
       (.I0(\processor/mem_exception ),
        .I1(\exception_context_out[ie1]_i_4_n_0 ),
        .I2(\exception_context_out[ie1]_i_6_n_0 ),
        .I3(\processor/mem_exception_context ),
        .I4(\processor/mem_csr_data [3]),
        .O(\processor/ex_exception_context ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \exception_context_out[ie1]_i_4 
       (.I0(\processor/mem_csr_address [4]),
        .I1(\processor/mem_csr_address [3]),
        .I2(\processor/mem_csr_address [7]),
        .I3(\processor/mem_csr_address [2]),
        .I4(\exception_context_out[ie1]_i_7_n_0 ),
        .I5(\exception_context_out[ie1]_i_8_n_0 ),
        .O(\exception_context_out[ie1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \exception_context_out[ie1]_i_5 
       (.I0(\processor/wb_exception_context[ie] ),
        .I1(\processor/wb_exception ),
        .I2(\processor/wb_csr_data [0]),
        .I3(\exception_context_out[ie1]_i_9_n_0 ),
        .I4(\processor/ie ),
        .O(\exception_context_out[ie1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \exception_context_out[ie1]_i_6 
       (.I0(\processor/wb_csr_data [3]),
        .I1(\exception_context_out[ie1]_i_9_n_0 ),
        .I2(\processor/ie1 ),
        .I3(\processor/wb_exception_context ),
        .I4(\processor/wb_exception ),
        .O(\exception_context_out[ie1]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0008)) 
    \exception_context_out[ie1]_i_7 
       (.I0(\processor/mem_csr_address [9]),
        .I1(\processor/mem_csr_address [8]),
        .I2(\processor/mem_csr_address [5]),
        .I3(\processor/mem_csr_address [6]),
        .O(\exception_context_out[ie1]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF1)) 
    \exception_context_out[ie1]_i_8 
       (.I0(\processor/mem_csr_write [1]),
        .I1(\processor/mem_csr_write [0]),
        .I2(\processor/mem_csr_address [0]),
        .I3(\processor/mem_csr_address [11]),
        .I4(\processor/mem_csr_address [1]),
        .I5(\processor/mem_csr_address [10]),
        .O(\exception_context_out[ie1]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \exception_context_out[ie1]_i_9 
       (.I0(\exception_context_out[ie1]_i_10_n_0 ),
        .I1(\exception_context_out[ie1]_i_11_n_0 ),
        .I2(\processor/wb_csr_address [2]),
        .O(\exception_context_out[ie1]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF000000FF00E2E2)) 
    \exception_context_out[ie]_i_1 
       (.I0(\processor/ex_exception_context[ie] ),
        .I1(\exception_context_out[ie]_i_2_n_0 ),
        .I2(\processor/ex_exception_context ),
        .I3(\processor/mem_exception_context[ie] ),
        .I4(reset),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(\exception_context_out[ie]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \exception_context_out[ie]_i_2 
       (.I0(\processor/ex_branch [2]),
        .I1(\processor/ex_branch [0]),
        .I2(\processor/ex_branch [1]),
        .O(\exception_context_out[ie]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABAA)) 
    exception_out_i_1
       (.I0(\mem_op[2]_i_5_n_0 ),
        .I1(\processor/ex_branch [1]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [2]),
        .O(\processor/memory/exception_out0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cache_hit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\icache/cache_hit0 ),
        .Q(\icache/cache_hit ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* IS_CLOCK_GATED *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* POWER_OPTED_CE = "ENBWREN=NEW" *) 
  (* RTL_RAM_BITS = "16384" *) 
  (* RTL_RAM_NAME = "cache_memory" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "511" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "71" *) 
  RAMB36E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .EN_ECC_READ("FALSE"),
    .EN_ECC_WRITE("FALSE"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(36'h000000000),
    .INIT_B(36'h000000000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_EXTENSION_A("NONE"),
    .RAM_EXTENSION_B("NONE"),
    .RAM_MODE("SDP"),
    .RDADDR_COLLISION_HWCONFIG("DELAYED_WRITE"),
    .READ_WIDTH_A(72),
    .READ_WIDTH_B(0),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(36'h000000000),
    .SRVAL_B(36'h000000000),
    .WRITE_MODE_A("READ_FIRST"),
    .WRITE_MODE_B("READ_FIRST"),
    .WRITE_WIDTH_A(0),
    .WRITE_WIDTH_B(72)) 
    \icache/cache_memory_reg_0 
       (.ADDRARDADDR({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,imem_address[10:4],\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .ADDRBWRADDR({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\icache/cl_load_address [10:4],\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CASCADEINA(\<const0>__0__0 ),
        .CASCADEINB(\<const0>__0__0 ),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI(\icache/load_buffer [31:0]),
        .DIBDI(\icache/load_buffer [63:32]),
        .DIPADIP(\icache/load_buffer [67:64]),
        .DIPBDIP(\icache/load_buffer [71:68]),
        .DOADO({\icache/current_cache_line [29:0],\icache/cache_memory_reg_0_n_51 ,\icache/cache_memory_reg_0_n_52 }),
        .DOBDO({\icache/current_cache_line [61:32],\icache/cache_memory_reg_0_n_83 ,\icache/cache_memory_reg_0_n_84 }),
        .DOPADOP({\icache/current_cache_line [65:64],\icache/cache_memory_reg_0_n_87 ,\icache/cache_memory_reg_0_n_88 }),
        .DOPBDOP(\icache/current_cache_line [69:66]),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\icache/store_cache_line_reg_n_0 ),
        .INJECTDBITERR(\<const0>__0__0 ),
        .INJECTSBITERR(\<const0>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\icache/store_cache_line_reg_n_0 ,\icache/store_cache_line_reg_n_0 ,\icache/store_cache_line_reg_n_0 ,\icache/store_cache_line_reg_n_0 ,\icache/store_cache_line_reg_n_0 ,\icache/store_cache_line_reg_n_0 ,\icache/store_cache_line_reg_n_0 ,\icache/store_cache_line_reg_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* IS_CLOCK_GATED *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* POWER_OPTED_CE = "ENBWREN=NEW" *) 
  (* RTL_RAM_BITS = "16384" *) 
  (* RTL_RAM_NAME = "cache_memory" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "511" *) 
  (* bram_slice_begin = "72" *) 
  (* bram_slice_end = "143" *) 
  RAMB36E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .EN_ECC_READ("FALSE"),
    .EN_ECC_WRITE("FALSE"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(36'h000000000),
    .INIT_B(36'h000000000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_EXTENSION_A("NONE"),
    .RAM_EXTENSION_B("NONE"),
    .RAM_MODE("SDP"),
    .RDADDR_COLLISION_HWCONFIG("DELAYED_WRITE"),
    .READ_WIDTH_A(72),
    .READ_WIDTH_B(0),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(36'h000000000),
    .SRVAL_B(36'h000000000),
    .WRITE_MODE_A("READ_FIRST"),
    .WRITE_MODE_B("READ_FIRST"),
    .WRITE_WIDTH_A(0),
    .WRITE_WIDTH_B(72)) 
    \icache/cache_memory_reg_1 
       (.ADDRARDADDR({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,imem_address[10:4],\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .ADDRBWRADDR({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\icache/cl_load_address [10:4],\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CASCADEINA(\<const0>__0__0 ),
        .CASCADEINB(\<const0>__0__0 ),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI(\icache/load_buffer [103:72]),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\icache/load_buffer [127:104]}),
        .DIPADIP({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\icache/current_cache_line [101:96],\icache/cache_memory_reg_1_n_27 ,\icache/cache_memory_reg_1_n_28 ,\icache/current_cache_line [93:70]}),
        .DOBDO({\icache/cache_memory_reg_1_n_53 ,\icache/cache_memory_reg_1_n_54 ,\icache/cache_memory_reg_1_n_55 ,\icache/cache_memory_reg_1_n_56 ,\icache/cache_memory_reg_1_n_57 ,\icache/cache_memory_reg_1_n_58 ,\icache/cache_memory_reg_1_n_59 ,\icache/cache_memory_reg_1_n_60 ,\icache/current_cache_line [125:102]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\icache/store_cache_line_reg_n_0 ),
        .INJECTDBITERR(\<const0>__0__0 ),
        .INJECTSBITERR(\<const0>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\icache/store_cache_line_reg_n_0 ,\icache/store_cache_line_reg_n_0 ,\icache/store_cache_line_reg_n_0 ,\icache/store_cache_line_reg_n_0 ,\icache/store_cache_line_reg_n_0 ,\icache/store_cache_line_reg_n_0 ,\icache/store_cache_line_reg_n_0 ,\icache/store_cache_line_reg_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_current_word_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(cl_current_word),
        .Q(\icache/cl_current_word_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_current_word_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\cl_current_word[1]_i_1_n_0 ),
        .Q(\icache/cl_current_word_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_current_word_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\cl_current_word[2]_i_1_n_0 ),
        .Q(\icache/cl_current_word_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[10] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[10]),
        .Q(\icache/cl_load_address [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[11] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[11]),
        .Q(\icache/cl_load_address [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[12] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[12]),
        .Q(\icache/cl_load_address [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[13] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[13]),
        .Q(\icache/cl_load_address [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[14] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[14]),
        .Q(\icache/cl_load_address [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[15] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[15]),
        .Q(\icache/cl_load_address [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[16] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[16]),
        .Q(\icache/cl_load_address [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[17] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[17]),
        .Q(\icache/cl_load_address [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[18] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[18]),
        .Q(\icache/cl_load_address [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[19] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[19]),
        .Q(\icache/cl_load_address [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[20] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[20]),
        .Q(\icache/cl_load_address [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[21] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[21]),
        .Q(\icache/cl_load_address [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[22] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[22]),
        .Q(\icache/cl_load_address [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[23] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[23]),
        .Q(\icache/cl_load_address [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[24] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[24]),
        .Q(\icache/cl_load_address [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[25] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[25]),
        .Q(\icache/cl_load_address [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[26] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[26]),
        .Q(\icache/cl_load_address [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[27] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[27]),
        .Q(\icache/cl_load_address [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[28] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[28]),
        .Q(\icache/cl_load_address [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[29] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[29]),
        .Q(\icache/cl_load_address [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[30] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[30]),
        .Q(\icache/cl_load_address [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[31] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[31]),
        .Q(\icache/cl_load_address [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[4] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[4]),
        .Q(\icache/cl_load_address [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[5] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[5]),
        .Q(\icache/cl_load_address [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[6] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[6]),
        .Q(\icache/cl_load_address [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[7] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[7]),
        .Q(\icache/cl_load_address [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[8] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[8]),
        .Q(\icache/cl_load_address [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/cl_load_address_reg[9] 
       (.C(clk),
        .CE(cl_load_address),
        .D(imem_address[9]),
        .Q(\icache/cl_load_address [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/input_address_word_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(imem_address[2]),
        .Q(\icache/input_address_word [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/input_address_word_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(imem_address[3]),
        .Q(\icache/input_address_word [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \icache/input_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\icache/input_carry_n_0 ,\icache/input_carry_n_1 ,\icache/input_carry_n_2 ,\icache/input_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({input_carry_i_1_n_0,input_carry_i_2_n_0,input_carry_i_3_n_0,input_carry_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \icache/input_carry__0 
       (.CI(\icache/input_carry_n_0 ),
        .CO({\icache/input_carry__0_n_0 ,\icache/to_std_logic ,\icache/input_carry__0_n_2 ,\icache/input_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const0>__0__0 ,input_carry__0_i_1_n_0,input_carry__0_i_2_n_0,input_carry__0_i_3_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[10]_i_1 
       (.I0(\icache/current_cache_line [104]),
        .I1(\icache/current_cache_line [40]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [72]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [8]),
        .O(imem_data[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[11]_i_1 
       (.I0(\icache/current_cache_line [105]),
        .I1(\icache/current_cache_line [41]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [73]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [9]),
        .O(imem_data[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[12]_i_1 
       (.I0(\icache/current_cache_line [106]),
        .I1(\icache/current_cache_line [42]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [74]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [10]),
        .O(imem_data[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[13]_i_1 
       (.I0(\icache/current_cache_line [107]),
        .I1(\icache/current_cache_line [43]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [75]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [11]),
        .O(imem_data[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[14]_i_1 
       (.I0(\icache/current_cache_line [108]),
        .I1(\icache/current_cache_line [44]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [76]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [12]),
        .O(imem_data[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[15]_i_1 
       (.I0(\icache/current_cache_line [109]),
        .I1(\icache/current_cache_line [45]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [77]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [13]),
        .O(imem_data[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[16]_i_1 
       (.I0(\icache/current_cache_line [110]),
        .I1(\icache/current_cache_line [46]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [78]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [14]),
        .O(imem_data[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[17]_i_1 
       (.I0(\icache/current_cache_line [111]),
        .I1(\icache/current_cache_line [47]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [79]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [15]),
        .O(imem_data[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[18]_i_1 
       (.I0(\icache/current_cache_line [112]),
        .I1(\icache/current_cache_line [48]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [80]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [16]),
        .O(imem_data[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[19]_i_1 
       (.I0(\icache/current_cache_line [113]),
        .I1(\icache/current_cache_line [49]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [81]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [17]),
        .O(imem_data[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[20]_i_1 
       (.I0(\icache/current_cache_line [114]),
        .I1(\icache/current_cache_line [50]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [82]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [18]),
        .O(imem_data[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[21]_i_1 
       (.I0(\icache/current_cache_line [115]),
        .I1(\icache/current_cache_line [51]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [83]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [19]),
        .O(imem_data[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[22]_i_1 
       (.I0(\icache/current_cache_line [116]),
        .I1(\icache/current_cache_line [52]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [84]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [20]),
        .O(imem_data[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[23]_i_1 
       (.I0(\icache/current_cache_line [117]),
        .I1(\icache/current_cache_line [53]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [85]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [21]),
        .O(imem_data[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[24]_i_1 
       (.I0(\icache/current_cache_line [118]),
        .I1(\icache/current_cache_line [54]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [86]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [22]),
        .O(imem_data[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[25]_i_1 
       (.I0(\icache/current_cache_line [119]),
        .I1(\icache/current_cache_line [55]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [87]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [23]),
        .O(imem_data[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[26]_i_1 
       (.I0(\icache/current_cache_line [120]),
        .I1(\icache/current_cache_line [56]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [88]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [24]),
        .O(imem_data[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[27]_i_1 
       (.I0(\icache/current_cache_line [121]),
        .I1(\icache/current_cache_line [57]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [89]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [25]),
        .O(imem_data[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[28]_i_1 
       (.I0(\icache/current_cache_line [122]),
        .I1(\icache/current_cache_line [58]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [90]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [26]),
        .O(imem_data[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[29]_i_1 
       (.I0(\icache/current_cache_line [123]),
        .I1(\icache/current_cache_line [59]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [91]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [27]),
        .O(imem_data[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[2]_i_1 
       (.I0(\icache/current_cache_line [96]),
        .I1(\icache/current_cache_line [32]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [64]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [0]),
        .O(imem_data[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[30]_i_1 
       (.I0(\icache/current_cache_line [124]),
        .I1(\icache/current_cache_line [60]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [92]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [28]),
        .O(imem_data[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[31]_i_2 
       (.I0(\icache/current_cache_line [125]),
        .I1(\icache/current_cache_line [61]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [93]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [29]),
        .O(imem_data[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[3]_i_1 
       (.I0(\icache/current_cache_line [97]),
        .I1(\icache/current_cache_line [33]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [65]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [1]),
        .O(imem_data[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[4]_i_1 
       (.I0(\icache/current_cache_line [98]),
        .I1(\icache/current_cache_line [34]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [66]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [2]),
        .O(imem_data[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[5]_i_1 
       (.I0(\icache/current_cache_line [99]),
        .I1(\icache/current_cache_line [35]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [67]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [3]),
        .O(imem_data[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[6]_i_1 
       (.I0(\icache/current_cache_line [100]),
        .I1(\icache/current_cache_line [36]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [68]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [4]),
        .O(imem_data[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[7]_i_1 
       (.I0(\icache/current_cache_line [101]),
        .I1(\icache/current_cache_line [37]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [69]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [5]),
        .O(imem_data[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[8]_i_1 
       (.I0(\icache/current_cache_line [102]),
        .I1(\icache/current_cache_line [38]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [70]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [6]),
        .O(imem_data[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \icache/instruction[9]_i_1 
       (.I0(\icache/current_cache_line [103]),
        .I1(\icache/current_cache_line [39]),
        .I2(\icache/input_address_word [0]),
        .I3(\icache/current_cache_line [71]),
        .I4(\icache/input_address_word [1]),
        .I5(\icache/current_cache_line [7]),
        .O(imem_data[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[0] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[64]_i_1_n_0 ),
        .Q(\icache/load_buffer [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[100] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(load_buffer),
        .Q(\icache/load_buffer [100]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[101] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[101]_i_1_n_0 ),
        .Q(\icache/load_buffer [101]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[102] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[102]_i_1_n_0 ),
        .Q(\icache/load_buffer [102]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[103] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[103]_i_1_n_0 ),
        .Q(\icache/load_buffer [103]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[104] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[104]_i_1_n_0 ),
        .Q(\icache/load_buffer [104]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[105] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[105]_i_1_n_0 ),
        .Q(\icache/load_buffer [105]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[106] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[106]_i_1_n_0 ),
        .Q(\icache/load_buffer [106]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[107] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[107]_i_1_n_0 ),
        .Q(\icache/load_buffer [107]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[108] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[108]_i_1_n_0 ),
        .Q(\icache/load_buffer [108]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[109] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[109]_i_1_n_0 ),
        .Q(\icache/load_buffer [109]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[10] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[74]_i_1_n_0 ),
        .Q(\icache/load_buffer [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[110] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[110]_i_1_n_0 ),
        .Q(\icache/load_buffer [110]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[111] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[111]_i_1_n_0 ),
        .Q(\icache/load_buffer [111]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[112] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[112]_i_1_n_0 ),
        .Q(\icache/load_buffer [112]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[113] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[113]_i_1_n_0 ),
        .Q(\icache/load_buffer [113]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[114] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[114]_i_1_n_0 ),
        .Q(\icache/load_buffer [114]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[115] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[115]_i_1_n_0 ),
        .Q(\icache/load_buffer [115]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[116] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[116]_i_1_n_0 ),
        .Q(\icache/load_buffer [116]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[117] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[117]_i_1_n_0 ),
        .Q(\icache/load_buffer [117]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[118] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[118]_i_1_n_0 ),
        .Q(\icache/load_buffer [118]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[119] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[119]_i_1_n_0 ),
        .Q(\icache/load_buffer [119]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[11] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[75]_i_1_n_0 ),
        .Q(\icache/load_buffer [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[120] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[120]_i_1_n_0 ),
        .Q(\icache/load_buffer [120]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[121] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[121]_i_1_n_0 ),
        .Q(\icache/load_buffer [121]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[122] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[122]_i_1_n_0 ),
        .Q(\icache/load_buffer [122]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[123] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[123]_i_1_n_0 ),
        .Q(\icache/load_buffer [123]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[124] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[124]_i_1_n_0 ),
        .Q(\icache/load_buffer [124]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[125] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[125]_i_1_n_0 ),
        .Q(\icache/load_buffer [125]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[126] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[126]_i_1_n_0 ),
        .Q(\icache/load_buffer [126]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[127] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[127]_i_2_n_0 ),
        .Q(\icache/load_buffer [127]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[12] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[76]_i_1_n_0 ),
        .Q(\icache/load_buffer [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[13] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[77]_i_1_n_0 ),
        .Q(\icache/load_buffer [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[14] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[78]_i_1_n_0 ),
        .Q(\icache/load_buffer [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[15] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[79]_i_1_n_0 ),
        .Q(\icache/load_buffer [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[16] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[80]_i_1_n_0 ),
        .Q(\icache/load_buffer [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[17] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[81]_i_1_n_0 ),
        .Q(\icache/load_buffer [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[18] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[82]_i_1_n_0 ),
        .Q(\icache/load_buffer [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[19] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[83]_i_1_n_0 ),
        .Q(\icache/load_buffer [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[1] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[65]_i_1_n_0 ),
        .Q(\icache/load_buffer [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[20] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[84]_i_1_n_0 ),
        .Q(\icache/load_buffer [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[21] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[85]_i_1_n_0 ),
        .Q(\icache/load_buffer [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[22] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[86]_i_1_n_0 ),
        .Q(\icache/load_buffer [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[23] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[87]_i_1_n_0 ),
        .Q(\icache/load_buffer [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[24] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[88]_i_1_n_0 ),
        .Q(\icache/load_buffer [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[25] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[89]_i_1_n_0 ),
        .Q(\icache/load_buffer [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[26] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[90]_i_1_n_0 ),
        .Q(\icache/load_buffer [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[27] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[91]_i_1_n_0 ),
        .Q(\icache/load_buffer [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[28] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[92]_i_1_n_0 ),
        .Q(\icache/load_buffer [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[29] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[93]_i_1_n_0 ),
        .Q(\icache/load_buffer [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[2] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[66]_i_1_n_0 ),
        .Q(\icache/load_buffer [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[30] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[94]_i_1_n_0 ),
        .Q(\icache/load_buffer [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[31] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[95]_i_2_n_0 ),
        .Q(\icache/load_buffer [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[32] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[96]_i_1_n_0 ),
        .Q(\icache/load_buffer [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[33] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[97]_i_1_n_0 ),
        .Q(\icache/load_buffer [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[34] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[98]_i_1_n_0 ),
        .Q(\icache/load_buffer [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[35] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[99]_i_1_n_0 ),
        .Q(\icache/load_buffer [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[36] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(load_buffer),
        .Q(\icache/load_buffer [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[37] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[101]_i_1_n_0 ),
        .Q(\icache/load_buffer [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[38] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[102]_i_1_n_0 ),
        .Q(\icache/load_buffer [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[39] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[103]_i_1_n_0 ),
        .Q(\icache/load_buffer [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[3] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[67]_i_1_n_0 ),
        .Q(\icache/load_buffer [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[40] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[104]_i_1_n_0 ),
        .Q(\icache/load_buffer [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[41] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[105]_i_1_n_0 ),
        .Q(\icache/load_buffer [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[42] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[106]_i_1_n_0 ),
        .Q(\icache/load_buffer [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[43] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[107]_i_1_n_0 ),
        .Q(\icache/load_buffer [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[44] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[108]_i_1_n_0 ),
        .Q(\icache/load_buffer [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[45] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[109]_i_1_n_0 ),
        .Q(\icache/load_buffer [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[46] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[110]_i_1_n_0 ),
        .Q(\icache/load_buffer [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[47] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[111]_i_1_n_0 ),
        .Q(\icache/load_buffer [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[48] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[112]_i_1_n_0 ),
        .Q(\icache/load_buffer [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[49] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[113]_i_1_n_0 ),
        .Q(\icache/load_buffer [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[4] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[68]_i_1_n_0 ),
        .Q(\icache/load_buffer [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[50] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[114]_i_1_n_0 ),
        .Q(\icache/load_buffer [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[51] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[115]_i_1_n_0 ),
        .Q(\icache/load_buffer [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[52] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[116]_i_1_n_0 ),
        .Q(\icache/load_buffer [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[53] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[117]_i_1_n_0 ),
        .Q(\icache/load_buffer [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[54] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[118]_i_1_n_0 ),
        .Q(\icache/load_buffer [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[55] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[119]_i_1_n_0 ),
        .Q(\icache/load_buffer [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[56] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[120]_i_1_n_0 ),
        .Q(\icache/load_buffer [56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[57] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[121]_i_1_n_0 ),
        .Q(\icache/load_buffer [57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[58] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[122]_i_1_n_0 ),
        .Q(\icache/load_buffer [58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[59] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[123]_i_1_n_0 ),
        .Q(\icache/load_buffer [59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[5] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[69]_i_1_n_0 ),
        .Q(\icache/load_buffer [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[60] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[124]_i_1_n_0 ),
        .Q(\icache/load_buffer [60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[61] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[125]_i_1_n_0 ),
        .Q(\icache/load_buffer [61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[62] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[126]_i_1_n_0 ),
        .Q(\icache/load_buffer [62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[63] 
       (.C(clk),
        .CE(\load_buffer[63]_i_1_n_0 ),
        .D(\load_buffer[127]_i_2_n_0 ),
        .Q(\icache/load_buffer [63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[64] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[64]_i_1_n_0 ),
        .Q(\icache/load_buffer [64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[65] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[65]_i_1_n_0 ),
        .Q(\icache/load_buffer [65]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[66] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[66]_i_1_n_0 ),
        .Q(\icache/load_buffer [66]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[67] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[67]_i_1_n_0 ),
        .Q(\icache/load_buffer [67]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[68] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[68]_i_1_n_0 ),
        .Q(\icache/load_buffer [68]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[69] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[69]_i_1_n_0 ),
        .Q(\icache/load_buffer [69]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[6] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[70]_i_1_n_0 ),
        .Q(\icache/load_buffer [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[70] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[70]_i_1_n_0 ),
        .Q(\icache/load_buffer [70]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[71] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[71]_i_1_n_0 ),
        .Q(\icache/load_buffer [71]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[72] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[72]_i_1_n_0 ),
        .Q(\icache/load_buffer [72]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[73] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[73]_i_1_n_0 ),
        .Q(\icache/load_buffer [73]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[74] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[74]_i_1_n_0 ),
        .Q(\icache/load_buffer [74]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[75] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[75]_i_1_n_0 ),
        .Q(\icache/load_buffer [75]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[76] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[76]_i_1_n_0 ),
        .Q(\icache/load_buffer [76]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[77] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[77]_i_1_n_0 ),
        .Q(\icache/load_buffer [77]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[78] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[78]_i_1_n_0 ),
        .Q(\icache/load_buffer [78]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[79] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[79]_i_1_n_0 ),
        .Q(\icache/load_buffer [79]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[7] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[71]_i_1_n_0 ),
        .Q(\icache/load_buffer [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[80] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[80]_i_1_n_0 ),
        .Q(\icache/load_buffer [80]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[81] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[81]_i_1_n_0 ),
        .Q(\icache/load_buffer [81]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[82] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[82]_i_1_n_0 ),
        .Q(\icache/load_buffer [82]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[83] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[83]_i_1_n_0 ),
        .Q(\icache/load_buffer [83]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[84] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[84]_i_1_n_0 ),
        .Q(\icache/load_buffer [84]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[85] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[85]_i_1_n_0 ),
        .Q(\icache/load_buffer [85]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[86] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[86]_i_1_n_0 ),
        .Q(\icache/load_buffer [86]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[87] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[87]_i_1_n_0 ),
        .Q(\icache/load_buffer [87]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[88] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[88]_i_1_n_0 ),
        .Q(\icache/load_buffer [88]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[89] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[89]_i_1_n_0 ),
        .Q(\icache/load_buffer [89]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[8] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[72]_i_1_n_0 ),
        .Q(\icache/load_buffer [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[90] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[90]_i_1_n_0 ),
        .Q(\icache/load_buffer [90]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[91] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[91]_i_1_n_0 ),
        .Q(\icache/load_buffer [91]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[92] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[92]_i_1_n_0 ),
        .Q(\icache/load_buffer [92]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[93] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[93]_i_1_n_0 ),
        .Q(\icache/load_buffer [93]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[94] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[94]_i_1_n_0 ),
        .Q(\icache/load_buffer [94]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[95] 
       (.C(clk),
        .CE(\load_buffer[95]_i_1_n_0 ),
        .D(\load_buffer[95]_i_2_n_0 ),
        .Q(\icache/load_buffer [95]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[96] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[96]_i_1_n_0 ),
        .Q(\icache/load_buffer [96]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[97] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[97]_i_1_n_0 ),
        .Q(\icache/load_buffer [97]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[98] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[98]_i_1_n_0 ),
        .Q(\icache/load_buffer [98]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[99] 
       (.C(clk),
        .CE(\load_buffer[127]_i_1_n_0 ),
        .D(\load_buffer[99]_i_1_n_0 ),
        .Q(\icache/load_buffer [99]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/load_buffer_reg[9] 
       (.C(clk),
        .CE(\load_buffer[31]_i_1_n_0 ),
        .D(\load_buffer[73]_i_1_n_0 ),
        .Q(\icache/load_buffer [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/read_ack_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(read_ack_i_1_n_0),
        .Q(\icache/read_ack ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/state_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(state),
        .Q(\icache/state_reg_n_0_ ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/state_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\state[1]_i_1_n_0 ),
        .Q(\icache/state_reg_n_0_[1] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/state_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\state[2]_i_1_n_0 ),
        .Q(\icache/state_reg_n_0_[2] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/store_cache_line_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(store_cache_line_i_1_n_0),
        .Q(\icache/store_cache_line_reg_n_0 ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \icache/tag_memory_reg_0_63_0_2 
       (.ADDRA(imem_address[9:4]),
        .ADDRB(imem_address[9:4]),
        .ADDRC(imem_address[9:4]),
        .ADDRD(\icache/cl_load_address [9:4]),
        .DIA(\icache/cl_load_address [11]),
        .DIB(\icache/cl_load_address [12]),
        .DIC(\icache/cl_load_address [13]),
        .DID(\<const0>__0__0 ),
        .DOA(\icache/tag_memory_reg_0_63_0_2_n_0 ),
        .DOB(\icache/tag_memory_reg_0_63_0_2_n_1 ),
        .DOC(\icache/tag_memory_reg_0_63_0_2_n_2 ),
        .WCLK(clk),
        .WE(tag_memory_reg_0_63_0_2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \icache/tag_memory_reg_0_63_12_14 
       (.ADDRA(imem_address[9:4]),
        .ADDRB(imem_address[9:4]),
        .ADDRC(imem_address[9:4]),
        .ADDRD(\icache/cl_load_address [9:4]),
        .DIA(\icache/cl_load_address [23]),
        .DIB(\icache/cl_load_address [24]),
        .DIC(\icache/cl_load_address [25]),
        .DID(\<const0>__0__0 ),
        .DOA(\icache/tag_memory_reg_0_63_12_14_n_0 ),
        .DOB(\icache/tag_memory_reg_0_63_12_14_n_1 ),
        .DOC(\icache/tag_memory_reg_0_63_12_14_n_2 ),
        .WCLK(clk),
        .WE(tag_memory_reg_0_63_0_2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \icache/tag_memory_reg_0_63_15_17 
       (.ADDRA(imem_address[9:4]),
        .ADDRB(imem_address[9:4]),
        .ADDRC(imem_address[9:4]),
        .ADDRD(\icache/cl_load_address [9:4]),
        .DIA(\icache/cl_load_address [26]),
        .DIB(\icache/cl_load_address [27]),
        .DIC(\icache/cl_load_address [28]),
        .DID(\<const0>__0__0 ),
        .DOA(\icache/tag_memory_reg_0_63_15_17_n_0 ),
        .DOB(\icache/tag_memory_reg_0_63_15_17_n_1 ),
        .DOC(\icache/tag_memory_reg_0_63_15_17_n_2 ),
        .WCLK(clk),
        .WE(tag_memory_reg_0_63_0_2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \icache/tag_memory_reg_0_63_18_20 
       (.ADDRA(imem_address[9:4]),
        .ADDRB(imem_address[9:4]),
        .ADDRC(imem_address[9:4]),
        .ADDRD(\icache/cl_load_address [9:4]),
        .DIA(\icache/cl_load_address [29]),
        .DIB(\icache/cl_load_address [30]),
        .DIC(\icache/cl_load_address [31]),
        .DID(\<const0>__0__0 ),
        .DOA(\icache/tag_memory_reg_0_63_18_20_n_0 ),
        .DOB(\icache/tag_memory_reg_0_63_18_20_n_1 ),
        .DOC(\icache/tag_memory_reg_0_63_18_20_n_2 ),
        .WCLK(clk),
        .WE(tag_memory_reg_0_63_0_2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \icache/tag_memory_reg_0_63_3_5 
       (.ADDRA(imem_address[9:4]),
        .ADDRB(imem_address[9:4]),
        .ADDRC(imem_address[9:4]),
        .ADDRD(\icache/cl_load_address [9:4]),
        .DIA(\icache/cl_load_address [14]),
        .DIB(\icache/cl_load_address [15]),
        .DIC(\icache/cl_load_address [16]),
        .DID(\<const0>__0__0 ),
        .DOA(\icache/tag_memory_reg_0_63_3_5_n_0 ),
        .DOB(\icache/tag_memory_reg_0_63_3_5_n_1 ),
        .DOC(\icache/tag_memory_reg_0_63_3_5_n_2 ),
        .WCLK(clk),
        .WE(tag_memory_reg_0_63_0_2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \icache/tag_memory_reg_0_63_6_8 
       (.ADDRA(imem_address[9:4]),
        .ADDRB(imem_address[9:4]),
        .ADDRC(imem_address[9:4]),
        .ADDRD(\icache/cl_load_address [9:4]),
        .DIA(\icache/cl_load_address [17]),
        .DIB(\icache/cl_load_address [18]),
        .DIC(\icache/cl_load_address [19]),
        .DID(\<const0>__0__0 ),
        .DOA(\icache/tag_memory_reg_0_63_6_8_n_0 ),
        .DOB(\icache/tag_memory_reg_0_63_6_8_n_1 ),
        .DOC(\icache/tag_memory_reg_0_63_6_8_n_2 ),
        .WCLK(clk),
        .WE(tag_memory_reg_0_63_0_2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \icache/tag_memory_reg_0_63_9_11 
       (.ADDRA(imem_address[9:4]),
        .ADDRB(imem_address[9:4]),
        .ADDRC(imem_address[9:4]),
        .ADDRD(\icache/cl_load_address [9:4]),
        .DIA(\icache/cl_load_address [20]),
        .DIB(\icache/cl_load_address [21]),
        .DIC(\icache/cl_load_address [22]),
        .DID(\<const0>__0__0 ),
        .DOA(\icache/tag_memory_reg_0_63_9_11_n_0 ),
        .DOB(\icache/tag_memory_reg_0_63_9_11_n_1 ),
        .DOC(\icache/tag_memory_reg_0_63_9_11_n_2 ),
        .WCLK(clk),
        .WE(tag_memory_reg_0_63_0_2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \icache/tag_memory_reg_64_127_0_2 
       (.ADDRA(imem_address[9:4]),
        .ADDRB(imem_address[9:4]),
        .ADDRC(imem_address[9:4]),
        .ADDRD(\icache/cl_load_address [9:4]),
        .DIA(\icache/cl_load_address [11]),
        .DIB(\icache/cl_load_address [12]),
        .DIC(\icache/cl_load_address [13]),
        .DID(\<const0>__0__0 ),
        .DOA(\icache/tag_memory_reg_64_127_0_2_n_0 ),
        .DOB(\icache/tag_memory_reg_64_127_0_2_n_1 ),
        .DOC(\icache/tag_memory_reg_64_127_0_2_n_2 ),
        .WCLK(clk),
        .WE(tag_memory_reg_64_127_0_2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \icache/tag_memory_reg_64_127_12_14 
       (.ADDRA(imem_address[9:4]),
        .ADDRB(imem_address[9:4]),
        .ADDRC(imem_address[9:4]),
        .ADDRD(\icache/cl_load_address [9:4]),
        .DIA(\icache/cl_load_address [23]),
        .DIB(\icache/cl_load_address [24]),
        .DIC(\icache/cl_load_address [25]),
        .DID(\<const0>__0__0 ),
        .DOA(\icache/tag_memory_reg_64_127_12_14_n_0 ),
        .DOB(\icache/tag_memory_reg_64_127_12_14_n_1 ),
        .DOC(\icache/tag_memory_reg_64_127_12_14_n_2 ),
        .WCLK(clk),
        .WE(tag_memory_reg_64_127_0_2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \icache/tag_memory_reg_64_127_15_17 
       (.ADDRA(imem_address[9:4]),
        .ADDRB(imem_address[9:4]),
        .ADDRC(imem_address[9:4]),
        .ADDRD(\icache/cl_load_address [9:4]),
        .DIA(\icache/cl_load_address [26]),
        .DIB(\icache/cl_load_address [27]),
        .DIC(\icache/cl_load_address [28]),
        .DID(\<const0>__0__0 ),
        .DOA(\icache/tag_memory_reg_64_127_15_17_n_0 ),
        .DOB(\icache/tag_memory_reg_64_127_15_17_n_1 ),
        .DOC(\icache/tag_memory_reg_64_127_15_17_n_2 ),
        .WCLK(clk),
        .WE(tag_memory_reg_64_127_0_2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \icache/tag_memory_reg_64_127_18_20 
       (.ADDRA(imem_address[9:4]),
        .ADDRB(imem_address[9:4]),
        .ADDRC(imem_address[9:4]),
        .ADDRD(\icache/cl_load_address [9:4]),
        .DIA(\icache/cl_load_address [29]),
        .DIB(\icache/cl_load_address [30]),
        .DIC(\icache/cl_load_address [31]),
        .DID(\<const0>__0__0 ),
        .DOA(\icache/tag_memory_reg_64_127_18_20_n_0 ),
        .DOB(\icache/tag_memory_reg_64_127_18_20_n_1 ),
        .DOC(\icache/tag_memory_reg_64_127_18_20_n_2 ),
        .WCLK(clk),
        .WE(tag_memory_reg_64_127_0_2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \icache/tag_memory_reg_64_127_3_5 
       (.ADDRA(imem_address[9:4]),
        .ADDRB(imem_address[9:4]),
        .ADDRC(imem_address[9:4]),
        .ADDRD(\icache/cl_load_address [9:4]),
        .DIA(\icache/cl_load_address [14]),
        .DIB(\icache/cl_load_address [15]),
        .DIC(\icache/cl_load_address [16]),
        .DID(\<const0>__0__0 ),
        .DOA(\icache/tag_memory_reg_64_127_3_5_n_0 ),
        .DOB(\icache/tag_memory_reg_64_127_3_5_n_1 ),
        .DOC(\icache/tag_memory_reg_64_127_3_5_n_2 ),
        .WCLK(clk),
        .WE(tag_memory_reg_64_127_0_2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \icache/tag_memory_reg_64_127_6_8 
       (.ADDRA(imem_address[9:4]),
        .ADDRB(imem_address[9:4]),
        .ADDRC(imem_address[9:4]),
        .ADDRD(\icache/cl_load_address [9:4]),
        .DIA(\icache/cl_load_address [17]),
        .DIB(\icache/cl_load_address [18]),
        .DIC(\icache/cl_load_address [19]),
        .DID(\<const0>__0__0 ),
        .DOA(\icache/tag_memory_reg_64_127_6_8_n_0 ),
        .DOB(\icache/tag_memory_reg_64_127_6_8_n_1 ),
        .DOC(\icache/tag_memory_reg_64_127_6_8_n_2 ),
        .WCLK(clk),
        .WE(tag_memory_reg_64_127_0_2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \icache/tag_memory_reg_64_127_9_11 
       (.ADDRA(imem_address[9:4]),
        .ADDRB(imem_address[9:4]),
        .ADDRC(imem_address[9:4]),
        .ADDRD(\icache/cl_load_address [9:4]),
        .DIA(\icache/cl_load_address [20]),
        .DIB(\icache/cl_load_address [21]),
        .DIC(\icache/cl_load_address [22]),
        .DID(\<const0>__0__0 ),
        .DOA(\icache/tag_memory_reg_64_127_9_11_n_0 ),
        .DOB(\icache/tag_memory_reg_64_127_9_11_n_1 ),
        .DOC(\icache/tag_memory_reg_64_127_9_11_n_2 ),
        .WCLK(clk),
        .WE(tag_memory_reg_64_127_0_2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(valid),
        .Q(\icache/valid [0]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[100] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[100]_i_1_n_0 ),
        .Q(\icache/valid [100]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[101] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[101]_i_1_n_0 ),
        .Q(\icache/valid [101]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[102] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[102]_i_1_n_0 ),
        .Q(\icache/valid [102]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[103] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[103]_i_1_n_0 ),
        .Q(\icache/valid [103]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[104] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[104]_i_1_n_0 ),
        .Q(\icache/valid [104]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[105] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[105]_i_1_n_0 ),
        .Q(\icache/valid [105]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[106] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[106]_i_1_n_0 ),
        .Q(\icache/valid [106]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[107] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[107]_i_1_n_0 ),
        .Q(\icache/valid [107]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[108] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[108]_i_1_n_0 ),
        .Q(\icache/valid [108]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[109] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[109]_i_1_n_0 ),
        .Q(\icache/valid [109]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[10]_i_1_n_0 ),
        .Q(\icache/valid [10]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[110] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[110]_i_1_n_0 ),
        .Q(\icache/valid [110]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[111] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[111]_i_1_n_0 ),
        .Q(\icache/valid [111]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[112] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[112]_i_1_n_0 ),
        .Q(\icache/valid [112]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[113] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[113]_i_1_n_0 ),
        .Q(\icache/valid [113]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[114] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[114]_i_1_n_0 ),
        .Q(\icache/valid [114]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[115] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[115]_i_1_n_0 ),
        .Q(\icache/valid [115]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[116] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[116]_i_1_n_0 ),
        .Q(\icache/valid [116]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[117] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[117]_i_1_n_0 ),
        .Q(\icache/valid [117]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[118] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[118]_i_1_n_0 ),
        .Q(\icache/valid [118]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[119] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[119]_i_1_n_0 ),
        .Q(\icache/valid [119]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[11]_i_1_n_0 ),
        .Q(\icache/valid [11]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[120] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[120]_i_1_n_0 ),
        .Q(\icache/valid [120]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[121] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[121]_i_1_n_0 ),
        .Q(\icache/valid [121]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[122] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[122]_i_1_n_0 ),
        .Q(\icache/valid [122]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[123] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[123]_i_1_n_0 ),
        .Q(\icache/valid [123]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[124] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[124]_i_1_n_0 ),
        .Q(\icache/valid [124]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[125] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[125]_i_1_n_0 ),
        .Q(\icache/valid [125]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[126] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[126]_i_1_n_0 ),
        .Q(\icache/valid [126]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[127] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[127]_i_1_n_0 ),
        .Q(\icache/valid [127]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[12]_i_1_n_0 ),
        .Q(\icache/valid [12]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[13]_i_1_n_0 ),
        .Q(\icache/valid [13]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[14]_i_1_n_0 ),
        .Q(\icache/valid [14]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[15]_i_1_n_0 ),
        .Q(\icache/valid [15]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[16]_i_1_n_0 ),
        .Q(\icache/valid [16]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[17]_i_1_n_0 ),
        .Q(\icache/valid [17]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[18]_i_1_n_0 ),
        .Q(\icache/valid [18]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[19]_i_1_n_0 ),
        .Q(\icache/valid [19]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[1]_i_1_n_0 ),
        .Q(\icache/valid [1]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[20]_i_1_n_0 ),
        .Q(\icache/valid [20]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[21]_i_1_n_0 ),
        .Q(\icache/valid [21]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[22]_i_1_n_0 ),
        .Q(\icache/valid [22]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[23]_i_1_n_0 ),
        .Q(\icache/valid [23]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[24]_i_1_n_0 ),
        .Q(\icache/valid [24]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[25]_i_1_n_0 ),
        .Q(\icache/valid [25]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[26]_i_1_n_0 ),
        .Q(\icache/valid [26]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[27]_i_1_n_0 ),
        .Q(\icache/valid [27]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[28]_i_1_n_0 ),
        .Q(\icache/valid [28]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[29]_i_1_n_0 ),
        .Q(\icache/valid [29]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[2]_i_1_n_0 ),
        .Q(\icache/valid [2]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[30]_i_1_n_0 ),
        .Q(\icache/valid [30]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[31]_i_1_n_0 ),
        .Q(\icache/valid [31]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[32]_i_1_n_0 ),
        .Q(\icache/valid [32]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[33]_i_1_n_0 ),
        .Q(\icache/valid [33]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[34]_i_1_n_0 ),
        .Q(\icache/valid [34]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[35]_i_1_n_0 ),
        .Q(\icache/valid [35]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[36]_i_1_n_0 ),
        .Q(\icache/valid [36]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[37]_i_1_n_0 ),
        .Q(\icache/valid [37]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[38]_i_1_n_0 ),
        .Q(\icache/valid [38]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[39]_i_1_n_0 ),
        .Q(\icache/valid [39]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[3]_i_1_n_0 ),
        .Q(\icache/valid [3]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[40]_i_1_n_0 ),
        .Q(\icache/valid [40]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[41]_i_1_n_0 ),
        .Q(\icache/valid [41]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[42]_i_1_n_0 ),
        .Q(\icache/valid [42]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[43]_i_1_n_0 ),
        .Q(\icache/valid [43]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[44]_i_1_n_0 ),
        .Q(\icache/valid [44]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[45]_i_1_n_0 ),
        .Q(\icache/valid [45]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[46]_i_1_n_0 ),
        .Q(\icache/valid [46]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[47]_i_1_n_0 ),
        .Q(\icache/valid [47]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[48]_i_1_n_0 ),
        .Q(\icache/valid [48]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[49]_i_1_n_0 ),
        .Q(\icache/valid [49]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[4]_i_1_n_0 ),
        .Q(\icache/valid [4]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[50]_i_1_n_0 ),
        .Q(\icache/valid [50]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[51]_i_1_n_0 ),
        .Q(\icache/valid [51]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[52]_i_1_n_0 ),
        .Q(\icache/valid [52]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[53]_i_1_n_0 ),
        .Q(\icache/valid [53]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[54]_i_1_n_0 ),
        .Q(\icache/valid [54]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[55]_i_1_n_0 ),
        .Q(\icache/valid [55]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[56]_i_1_n_0 ),
        .Q(\icache/valid [56]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[57]_i_1_n_0 ),
        .Q(\icache/valid [57]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[58]_i_1_n_0 ),
        .Q(\icache/valid [58]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[59]_i_1_n_0 ),
        .Q(\icache/valid [59]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[5]_i_1_n_0 ),
        .Q(\icache/valid [5]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[60]_i_1_n_0 ),
        .Q(\icache/valid [60]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[61]_i_1_n_0 ),
        .Q(\icache/valid [61]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[62]_i_1_n_0 ),
        .Q(\icache/valid [62]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[63]_i_1_n_0 ),
        .Q(\icache/valid [63]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[64] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[64]_i_1_n_0 ),
        .Q(\icache/valid [64]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[65] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[65]_i_1_n_0 ),
        .Q(\icache/valid [65]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[66] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[66]_i_1_n_0 ),
        .Q(\icache/valid [66]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[67] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[67]_i_1_n_0 ),
        .Q(\icache/valid [67]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[68] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[68]_i_1_n_0 ),
        .Q(\icache/valid [68]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[69] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[69]_i_1_n_0 ),
        .Q(\icache/valid [69]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[6]_i_1_n_0 ),
        .Q(\icache/valid [6]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[70] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[70]_i_1_n_0 ),
        .Q(\icache/valid [70]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[71] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[71]_i_1_n_0 ),
        .Q(\icache/valid [71]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[72] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[72]_i_1_n_0 ),
        .Q(\icache/valid [72]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[73] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[73]_i_1_n_0 ),
        .Q(\icache/valid [73]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[74] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[74]_i_1_n_0 ),
        .Q(\icache/valid [74]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[75] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[75]_i_1_n_0 ),
        .Q(\icache/valid [75]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[76] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[76]_i_1_n_0 ),
        .Q(\icache/valid [76]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[77] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[77]_i_1_n_0 ),
        .Q(\icache/valid [77]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[78] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[78]_i_1_n_0 ),
        .Q(\icache/valid [78]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[79] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[79]_i_1_n_0 ),
        .Q(\icache/valid [79]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[7]_i_1_n_0 ),
        .Q(\icache/valid [7]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[80] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[80]_i_1_n_0 ),
        .Q(\icache/valid [80]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[81] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[81]_i_1_n_0 ),
        .Q(\icache/valid [81]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[82] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[82]_i_1_n_0 ),
        .Q(\icache/valid [82]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[83] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[83]_i_1_n_0 ),
        .Q(\icache/valid [83]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[84] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[84]_i_1_n_0 ),
        .Q(\icache/valid [84]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[85] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[85]_i_1_n_0 ),
        .Q(\icache/valid [85]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[86] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[86]_i_1_n_0 ),
        .Q(\icache/valid [86]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[87] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[87]_i_1_n_0 ),
        .Q(\icache/valid [87]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[88] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[88]_i_1_n_0 ),
        .Q(\icache/valid [88]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[89] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[89]_i_1_n_0 ),
        .Q(\icache/valid [89]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[8]_i_1_n_0 ),
        .Q(\icache/valid [8]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[90] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[90]_i_1_n_0 ),
        .Q(\icache/valid [90]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[91] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[91]_i_1_n_0 ),
        .Q(\icache/valid [91]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[92] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[92]_i_1_n_0 ),
        .Q(\icache/valid [92]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[93] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[93]_i_1_n_0 ),
        .Q(\icache/valid [93]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[94] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[94]_i_1_n_0 ),
        .Q(\icache/valid [94]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[95] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[95]_i_1_n_0 ),
        .Q(\icache/valid [95]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[96] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[96]_i_1_n_0 ),
        .Q(\icache/valid [96]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[97] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[97]_i_1_n_0 ),
        .Q(\icache/valid [97]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[98] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[98]_i_1_n_0 ),
        .Q(\icache/valid [98]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[99] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[99]_i_1_n_0 ),
        .Q(\icache/valid [99]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/valid_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\valid[9]_i_1_n_0 ),
        .Q(\icache/valid [9]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][10] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(wb_outputs),
        .Q(\icache_outputs[adr] [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][11] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][11]_i_1_n_0 ),
        .Q(\icache_outputs[adr] [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][12] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][12]_i_1__0_n_0 ),
        .Q(\icache_outputs[adr] [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][13] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][13]_i_1__0_n_0 ),
        .Q(\icache_outputs[adr] [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][14] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][14]_i_1_n_0 ),
        .Q(\icache_outputs[adr] [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][15] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][15]_i_1__0_n_0 ),
        .Q(\icache_outputs[adr] [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][16] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][16]_i_1__0_n_0 ),
        .Q(\icache_outputs[adr] [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][17] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][17]_i_1_n_0 ),
        .Q(\icache_outputs[adr] [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][18] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][18]_i_1__0_n_0 ),
        .Q(\icache_outputs[adr] [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][19] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][19]_i_1__0_n_0 ),
        .Q(\icache_outputs[adr] [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][20] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][20]_i_1_n_0 ),
        .Q(\icache_outputs[adr] [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][21] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][21]_i_1__0_n_0 ),
        .Q(\icache_outputs[adr] [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][22] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][22]_i_1__0_n_0 ),
        .Q(\icache_outputs[adr] [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][23] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][23]_i_1_n_0 ),
        .Q(\icache_outputs[adr] [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][24] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][24]_i_1__0_n_0 ),
        .Q(\icache_outputs[adr] [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][25] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][25]_i_1__0_n_0 ),
        .Q(\icache_outputs[adr] [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][26] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][26]_i_1_n_0 ),
        .Q(\icache_outputs[adr] [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][27] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][27]_i_1__0_n_0 ),
        .Q(\icache_outputs[adr] [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][28] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][28]_i_1__0_n_0 ),
        .Q(\icache_outputs[adr] [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][29] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][29]_i_1_n_0 ),
        .Q(\icache_outputs[adr] [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][2] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][2]_i_1__0_n_0 ),
        .Q(\icache_outputs[adr] [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][30] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][30]_i_1__0_n_0 ),
        .Q(\icache_outputs[adr] [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][31] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][31]_i_2__0_n_0 ),
        .Q(\icache_outputs[adr] [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][3] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][3]_i_1__0_n_0 ),
        .Q(\icache_outputs[adr] [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][4] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][4]_i_1_n_0 ),
        .Q(\icache_outputs[adr] [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][5] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][5]_i_1_n_0 ),
        .Q(\icache_outputs[adr] [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][6] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][6]_i_1__0_n_0 ),
        .Q(\icache_outputs[adr] [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][7] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][7]_i_1__0_n_0 ),
        .Q(\icache_outputs[adr] [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][8] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][8]_i_1_n_0 ),
        .Q(\icache_outputs[adr] [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[adr][9] 
       (.C(clk),
        .CE(\wb_outputs[adr][31]_i_1__0_n_0 ),
        .D(\wb_outputs[adr][9]_i_1_n_0 ),
        .Q(\icache_outputs[adr] [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[cyc] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\wb_outputs[cyc]_i_1__0_n_0 ),
        .Q(icache_outputs),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[sel][3] 
       (.C(clk),
        .CE(cl_load_address),
        .D(\icache/p_1_in10_out ),
        .Q(\icache_outputs[sel] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \icache/wb_outputs_reg[stb] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\wb_outputs[stb]_i_1_n_0 ),
        .Q(\icache_outputs[stb] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFB08FFFFFB080000)) 
    ie1_i_1
       (.I0(\processor/csr_unit/ie1__0 ),
        .I1(\processor/csr_unit/tohost_data1__0 ),
        .I2(\mtime_compare[31]_i_3_n_0 ),
        .I3(\processor/wb_exception_context ),
        .I4(ie_i_3_n_0),
        .I5(\processor/ie1 ),
        .O(ie1_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00FF01FF00FE00)) 
    ie1_i_2
       (.I0(\processor/wb_csr_address [4]),
        .I1(\processor/wb_csr_address [1]),
        .I2(\processor/wb_csr_address [3]),
        .I3(\processor/wb_exception_context ),
        .I4(\processor/wb_csr_address [5]),
        .I5(ie1_i_3_n_0),
        .O(\processor/csr_unit/ie1__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF0F1F0E0)) 
    ie1_i_3
       (.I0(\processor/wb_csr_address [2]),
        .I1(\processor/wb_csr_address [6]),
        .I2(\processor/wb_exception_context ),
        .I3(\processor/wb_csr_address [0]),
        .I4(\processor/wb_csr_data [3]),
        .O(ie1_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFB08FFFFFB080000)) 
    ie_i_1
       (.I0(\processor/csr_unit/ie__7 ),
        .I1(\processor/csr_unit/tohost_data1__0 ),
        .I2(\mtime_compare[31]_i_3_n_0 ),
        .I3(\processor/wb_exception_context[ie] ),
        .I4(ie_i_3_n_0),
        .I5(\processor/ie ),
        .O(ie_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00FF01FF00FE00)) 
    ie_i_2
       (.I0(\processor/wb_csr_address [4]),
        .I1(\processor/wb_csr_address [1]),
        .I2(\processor/wb_csr_address [3]),
        .I3(\processor/wb_exception_context[ie] ),
        .I4(\processor/wb_csr_address [5]),
        .I5(ie_i_4_n_0),
        .O(\processor/csr_unit/ie__7 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00010000)) 
    ie_i_3
       (.I0(ie_i_5_n_0),
        .I1(\processor/wb_csr_address [5]),
        .I2(\processor/wb_csr_address [4]),
        .I3(\processor/wb_csr_address [6]),
        .I4(ie_i_6_n_0),
        .I5(\processor/wb_exception ),
        .O(ie_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF0F1F0E0)) 
    ie_i_4
       (.I0(\processor/wb_csr_address [2]),
        .I1(\processor/wb_csr_address [6]),
        .I2(\processor/wb_exception_context[ie] ),
        .I3(\processor/wb_csr_address [0]),
        .I4(\processor/wb_csr_data [0]),
        .O(ie_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    ie_i_5
       (.I0(\processor/wb_csr_address [2]),
        .I1(\processor/wb_csr_address [3]),
        .I2(\processor/wb_csr_address [0]),
        .I3(\processor/wb_csr_address [1]),
        .O(ie_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    ie_i_6
       (.I0(\processor/csr_unit/tohost_data1__0 ),
        .I1(\processor/wb_csr_address [8]),
        .I2(\processor/wb_csr_address [7]),
        .I3(\processor/wb_csr_address [10]),
        .I4(\processor/wb_csr_address [11]),
        .I5(\processor/wb_csr_address [9]),
        .O(ie_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4004400405040004)) 
    \immediate[0]_i_2 
       (.I0(\processor/decode/instruction_reg_n_0_[3] ),
        .I1(\processor/id_shamt [0]),
        .I2(\processor/decode/instruction_reg_n_0_[6] ),
        .I3(\processor/decode/instruction_reg_n_0_[5] ),
        .I4(\processor/id_rd_address [0]),
        .I5(\processor/decode/instruction_reg_n_0_[4] ),
        .O(immediate));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h10000000)) 
    \immediate[0]_i_3 
       (.I0(\processor/decode/instruction_reg_n_0_[4] ),
        .I1(\processor/decode/instruction_reg_n_0_[3] ),
        .I2(\processor/decode/instruction_reg_n_0_[5] ),
        .I3(\processor/decode/instruction_reg_n_0_[6] ),
        .I4(\processor/id_shamt [0]),
        .O(\immediate[0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8AAA8AAAAAAA0A80)) 
    \immediate[10]_i_1 
       (.I0(\mem_size[1]_i_1_n_0 ),
        .I1(\processor/decode/instruction_reg_n_0_[4] ),
        .I2(\processor/decode/instruction_reg_n_0_[5] ),
        .I3(\processor/decode/instruction_reg_n_0_[6] ),
        .I4(\processor/decode/instruction_reg_n_0_[3] ),
        .I5(\processor/decode/instruction_reg_n_0_ ),
        .O(\immediate[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000008484E444)) 
    \immediate[11]_i_2 
       (.I0(\processor/decode/instruction_reg_n_0_[6] ),
        .I1(data0[31]),
        .I2(\processor/decode/instruction_reg_n_0_[5] ),
        .I3(\processor/id_rd_address [0]),
        .I4(\processor/decode/instruction_reg_n_0_[4] ),
        .I5(\processor/decode/instruction_reg_n_0_[3] ),
        .O(\immediate[11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0808080000000800)) 
    \immediate[11]_i_3 
       (.I0(\processor/decode/instruction_reg_n_0_[5] ),
        .I1(\processor/decode/instruction_reg_n_0_[6] ),
        .I2(\processor/decode/instruction_reg_n_0_[4] ),
        .I3(data0[31]),
        .I4(\processor/decode/instruction_reg_n_0_[3] ),
        .I5(\processor/id_shamt [0]),
        .O(\immediate[11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4A404540AF000500)) 
    \immediate[12]_i_2 
       (.I0(\processor/decode/instruction_reg_n_0_[6] ),
        .I1(\processor/id_funct3 [0]),
        .I2(\processor/decode/instruction_reg_n_0_ ),
        .I3(data0[31]),
        .I4(\processor/decode/instruction_reg_n_0_[5] ),
        .I5(\processor/decode/instruction_reg_n_0_[4] ),
        .O(\immediate[12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h40000000)) 
    \immediate[12]_i_3 
       (.I0(\processor/decode/instruction_reg_n_0_[4] ),
        .I1(\processor/id_funct3 [0]),
        .I2(\processor/decode/instruction_reg_n_0_ ),
        .I3(\processor/decode/instruction_reg_n_0_[6] ),
        .I4(\processor/decode/instruction_reg_n_0_[5] ),
        .O(\immediate[12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4A404540AF000500)) 
    \immediate[13]_i_2 
       (.I0(\processor/decode/instruction_reg_n_0_[6] ),
        .I1(\processor/id_funct3 [1]),
        .I2(\processor/decode/instruction_reg_n_0_ ),
        .I3(data0[31]),
        .I4(\processor/decode/instruction_reg_n_0_[5] ),
        .I5(\processor/decode/instruction_reg_n_0_[4] ),
        .O(\immediate[13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h40000000)) 
    \immediate[13]_i_3 
       (.I0(\processor/decode/instruction_reg_n_0_[4] ),
        .I1(\processor/id_funct3 [1]),
        .I2(\processor/decode/instruction_reg_n_0_ ),
        .I3(\processor/decode/instruction_reg_n_0_[6] ),
        .I4(\processor/decode/instruction_reg_n_0_[5] ),
        .O(\immediate[13]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4A404540AF000500)) 
    \immediate[14]_i_2 
       (.I0(\processor/decode/instruction_reg_n_0_[6] ),
        .I1(\processor/id_csr_use_immediate ),
        .I2(\processor/decode/instruction_reg_n_0_ ),
        .I3(data0[31]),
        .I4(\processor/decode/instruction_reg_n_0_[5] ),
        .I5(\processor/decode/instruction_reg_n_0_[4] ),
        .O(\immediate[14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h40000000)) 
    \immediate[14]_i_3 
       (.I0(\processor/decode/instruction_reg_n_0_[4] ),
        .I1(\processor/id_csr_use_immediate ),
        .I2(\processor/decode/instruction_reg_n_0_ ),
        .I3(\processor/decode/instruction_reg_n_0_[6] ),
        .I4(\processor/decode/instruction_reg_n_0_[5] ),
        .O(\immediate[14]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4A404540AF000500)) 
    \immediate[15]_i_2 
       (.I0(\processor/decode/instruction_reg_n_0_[6] ),
        .I1(\processor/id_rs1_address [0]),
        .I2(\processor/decode/instruction_reg_n_0_ ),
        .I3(data0[31]),
        .I4(\processor/decode/instruction_reg_n_0_[5] ),
        .I5(\processor/decode/instruction_reg_n_0_[4] ),
        .O(\immediate[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h40000000)) 
    \immediate[15]_i_3 
       (.I0(\processor/decode/instruction_reg_n_0_[4] ),
        .I1(\processor/id_rs1_address [0]),
        .I2(\processor/decode/instruction_reg_n_0_ ),
        .I3(\processor/decode/instruction_reg_n_0_[6] ),
        .I4(\processor/decode/instruction_reg_n_0_[5] ),
        .O(\immediate[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4A404540AF000500)) 
    \immediate[16]_i_2 
       (.I0(\processor/decode/instruction_reg_n_0_[6] ),
        .I1(\processor/id_rs1_address [1]),
        .I2(\processor/decode/instruction_reg_n_0_ ),
        .I3(data0[31]),
        .I4(\processor/decode/instruction_reg_n_0_[5] ),
        .I5(\processor/decode/instruction_reg_n_0_[4] ),
        .O(\immediate[16]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h40000000)) 
    \immediate[16]_i_3 
       (.I0(\processor/decode/instruction_reg_n_0_[4] ),
        .I1(\processor/id_rs1_address [1]),
        .I2(\processor/decode/instruction_reg_n_0_ ),
        .I3(\processor/decode/instruction_reg_n_0_[6] ),
        .I4(\processor/decode/instruction_reg_n_0_[5] ),
        .O(\immediate[16]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4A404540AF000500)) 
    \immediate[17]_i_2 
       (.I0(\processor/decode/instruction_reg_n_0_[6] ),
        .I1(\processor/id_rs1_address [2]),
        .I2(\processor/decode/instruction_reg_n_0_ ),
        .I3(data0[31]),
        .I4(\processor/decode/instruction_reg_n_0_[5] ),
        .I5(\processor/decode/instruction_reg_n_0_[4] ),
        .O(\immediate[17]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h40000000)) 
    \immediate[17]_i_3 
       (.I0(\processor/decode/instruction_reg_n_0_[4] ),
        .I1(\processor/id_rs1_address [2]),
        .I2(\processor/decode/instruction_reg_n_0_ ),
        .I3(\processor/decode/instruction_reg_n_0_[6] ),
        .I4(\processor/decode/instruction_reg_n_0_[5] ),
        .O(\immediate[17]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4A404540AF000500)) 
    \immediate[18]_i_2 
       (.I0(\processor/decode/instruction_reg_n_0_[6] ),
        .I1(\processor/id_rs1_address [3]),
        .I2(\processor/decode/instruction_reg_n_0_ ),
        .I3(data0[31]),
        .I4(\processor/decode/instruction_reg_n_0_[5] ),
        .I5(\processor/decode/instruction_reg_n_0_[4] ),
        .O(\immediate[18]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h40000000)) 
    \immediate[18]_i_3 
       (.I0(\processor/decode/instruction_reg_n_0_[4] ),
        .I1(\processor/id_rs1_address [3]),
        .I2(\processor/decode/instruction_reg_n_0_ ),
        .I3(\processor/decode/instruction_reg_n_0_[6] ),
        .I4(\processor/decode/instruction_reg_n_0_[5] ),
        .O(\immediate[18]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4A404540AF000500)) 
    \immediate[19]_i_2 
       (.I0(\processor/decode/instruction_reg_n_0_[6] ),
        .I1(\processor/id_rs1_address [4]),
        .I2(\processor/decode/instruction_reg_n_0_ ),
        .I3(data0[31]),
        .I4(\processor/decode/instruction_reg_n_0_[5] ),
        .I5(\processor/decode/instruction_reg_n_0_[4] ),
        .O(\immediate[19]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h40000000)) 
    \immediate[19]_i_3 
       (.I0(\processor/decode/instruction_reg_n_0_[4] ),
        .I1(\processor/id_rs1_address [4]),
        .I2(\processor/decode/instruction_reg_n_0_ ),
        .I3(\processor/decode/instruction_reg_n_0_[6] ),
        .I4(\processor/decode/instruction_reg_n_0_[5] ),
        .O(\immediate[19]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4000FFFF40000000)) 
    \immediate[1]_i_1 
       (.I0(\processor/decode/instruction_reg_n_0_[4] ),
        .I1(\processor/decode/instruction_reg_n_0_[6] ),
        .I2(\processor/id_shamt [1]),
        .I3(\processor/decode/instruction_reg_n_0_[5] ),
        .I4(\processor/decode/instruction_reg_n_0_ ),
        .I5(\immediate[1]_i_2_n_0 ),
        .O(\processor/id_immediate [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000008484F404)) 
    \immediate[1]_i_2 
       (.I0(\processor/decode/instruction_reg_n_0_[6] ),
        .I1(\processor/id_shamt [1]),
        .I2(\processor/decode/instruction_reg_n_0_[5] ),
        .I3(\processor/id_rd_address [1]),
        .I4(\processor/decode/instruction_reg_n_0_[4] ),
        .I5(\processor/decode/instruction_reg_n_0_[3] ),
        .O(\immediate[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2F20FFFF2F200000)) 
    \immediate[20]_i_1 
       (.I0(\processor/id_shamt [0]),
        .I1(\immediate[30]_i_2_n_0 ),
        .I2(\processor/decode/instruction_reg_n_0_[4] ),
        .I3(\immediate[30]_i_3_n_0 ),
        .I4(\processor/decode/instruction_reg_n_0_ ),
        .I5(\immediate[30]_i_4_n_0 ),
        .O(\processor/id_immediate [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2F20FFFF2F200000)) 
    \immediate[21]_i_1 
       (.I0(\processor/id_shamt [1]),
        .I1(\immediate[30]_i_2_n_0 ),
        .I2(\processor/decode/instruction_reg_n_0_[4] ),
        .I3(\immediate[30]_i_3_n_0 ),
        .I4(\processor/decode/instruction_reg_n_0_ ),
        .I5(\immediate[30]_i_4_n_0 ),
        .O(\processor/id_immediate [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2F20FFFF2F200000)) 
    \immediate[22]_i_1 
       (.I0(\processor/id_shamt [2]),
        .I1(\immediate[30]_i_2_n_0 ),
        .I2(\processor/decode/instruction_reg_n_0_[4] ),
        .I3(\immediate[30]_i_3_n_0 ),
        .I4(\processor/decode/instruction_reg_n_0_ ),
        .I5(\immediate[30]_i_4_n_0 ),
        .O(\processor/id_immediate [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2F20FFFF2F200000)) 
    \immediate[23]_i_1 
       (.I0(\processor/id_shamt [3]),
        .I1(\immediate[30]_i_2_n_0 ),
        .I2(\processor/decode/instruction_reg_n_0_[4] ),
        .I3(\immediate[30]_i_3_n_0 ),
        .I4(\processor/decode/instruction_reg_n_0_ ),
        .I5(\immediate[30]_i_4_n_0 ),
        .O(\processor/id_immediate [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2F20FFFF2F200000)) 
    \immediate[24]_i_1 
       (.I0(\processor/id_shamt [4]),
        .I1(\immediate[30]_i_2_n_0 ),
        .I2(\processor/decode/instruction_reg_n_0_[4] ),
        .I3(\immediate[30]_i_3_n_0 ),
        .I4(\processor/decode/instruction_reg_n_0_ ),
        .I5(\immediate[30]_i_4_n_0 ),
        .O(\processor/id_immediate [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2F20FFFF2F200000)) 
    \immediate[25]_i_1 
       (.I0(data0[25]),
        .I1(\immediate[30]_i_2_n_0 ),
        .I2(\processor/decode/instruction_reg_n_0_[4] ),
        .I3(\immediate[30]_i_3_n_0 ),
        .I4(\processor/decode/instruction_reg_n_0_ ),
        .I5(\immediate[30]_i_4_n_0 ),
        .O(\processor/id_immediate [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2F20FFFF2F200000)) 
    \immediate[26]_i_1 
       (.I0(data0[26]),
        .I1(\immediate[30]_i_2_n_0 ),
        .I2(\processor/decode/instruction_reg_n_0_[4] ),
        .I3(\immediate[30]_i_3_n_0 ),
        .I4(\processor/decode/instruction_reg_n_0_ ),
        .I5(\immediate[30]_i_4_n_0 ),
        .O(\processor/id_immediate [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2F20FFFF2F200000)) 
    \immediate[27]_i_1 
       (.I0(data0[27]),
        .I1(\immediate[30]_i_2_n_0 ),
        .I2(\processor/decode/instruction_reg_n_0_[4] ),
        .I3(\immediate[30]_i_3_n_0 ),
        .I4(\processor/decode/instruction_reg_n_0_ ),
        .I5(\immediate[30]_i_4_n_0 ),
        .O(\processor/id_immediate [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2F20FFFF2F200000)) 
    \immediate[28]_i_1 
       (.I0(data0[28]),
        .I1(\immediate[30]_i_2_n_0 ),
        .I2(\processor/decode/instruction_reg_n_0_[4] ),
        .I3(\immediate[30]_i_3_n_0 ),
        .I4(\processor/decode/instruction_reg_n_0_ ),
        .I5(\immediate[30]_i_4_n_0 ),
        .O(\processor/id_immediate [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2F20FFFF2F200000)) 
    \immediate[29]_i_1 
       (.I0(data0[29]),
        .I1(\immediate[30]_i_2_n_0 ),
        .I2(\processor/decode/instruction_reg_n_0_[4] ),
        .I3(\immediate[30]_i_3_n_0 ),
        .I4(\processor/decode/instruction_reg_n_0_ ),
        .I5(\immediate[30]_i_4_n_0 ),
        .O(\processor/id_immediate [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4000FFFF40000000)) 
    \immediate[2]_i_1 
       (.I0(\processor/decode/instruction_reg_n_0_[4] ),
        .I1(\processor/decode/instruction_reg_n_0_[6] ),
        .I2(\processor/id_shamt [2]),
        .I3(\processor/decode/instruction_reg_n_0_[5] ),
        .I4(\processor/decode/instruction_reg_n_0_ ),
        .I5(\immediate[2]_i_2_n_0 ),
        .O(\processor/id_immediate [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000008484F404)) 
    \immediate[2]_i_2 
       (.I0(\processor/decode/instruction_reg_n_0_[6] ),
        .I1(\processor/id_shamt [2]),
        .I2(\processor/decode/instruction_reg_n_0_[5] ),
        .I3(\processor/id_rd_address [2]),
        .I4(\processor/decode/instruction_reg_n_0_[4] ),
        .I5(\processor/decode/instruction_reg_n_0_[3] ),
        .O(\immediate[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2F20FFFF2F200000)) 
    \immediate[30]_i_1 
       (.I0(data0[30]),
        .I1(\immediate[30]_i_2_n_0 ),
        .I2(\processor/decode/instruction_reg_n_0_[4] ),
        .I3(\immediate[30]_i_3_n_0 ),
        .I4(\processor/decode/instruction_reg_n_0_ ),
        .I5(\immediate[30]_i_4_n_0 ),
        .O(\processor/id_immediate [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \immediate[30]_i_2 
       (.I0(\processor/decode/instruction_reg_n_0_[6] ),
        .I1(\processor/decode/instruction_reg_n_0_[3] ),
        .O(\immediate[30]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \immediate[30]_i_3 
       (.I0(\processor/decode/instruction_reg_n_0_[6] ),
        .I1(\processor/decode/instruction_reg_n_0_[5] ),
        .I2(data0[31]),
        .O(\immediate[30]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h20220202)) 
    \immediate[30]_i_4 
       (.I0(data0[31]),
        .I1(\processor/decode/instruction_reg_n_0_[3] ),
        .I2(\processor/decode/instruction_reg_n_0_[6] ),
        .I3(\processor/decode/instruction_reg_n_0_[4] ),
        .I4(\processor/decode/instruction_reg_n_0_[5] ),
        .O(\immediate[30]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04088C04000C0004)) 
    \immediate[31]_i_1 
       (.I0(\processor/decode/instruction_reg_n_0_ ),
        .I1(data0[31]),
        .I2(\processor/decode/instruction_reg_n_0_[3] ),
        .I3(\processor/decode/instruction_reg_n_0_[6] ),
        .I4(\processor/decode/instruction_reg_n_0_[4] ),
        .I5(\processor/decode/instruction_reg_n_0_[5] ),
        .O(\processor/id_immediate [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4000FFFF40000000)) 
    \immediate[3]_i_1 
       (.I0(\processor/decode/instruction_reg_n_0_[4] ),
        .I1(\processor/decode/instruction_reg_n_0_[6] ),
        .I2(\processor/id_shamt [3]),
        .I3(\processor/decode/instruction_reg_n_0_[5] ),
        .I4(\processor/decode/instruction_reg_n_0_ ),
        .I5(\immediate[3]_i_2_n_0 ),
        .O(\processor/id_immediate [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000008484F404)) 
    \immediate[3]_i_2 
       (.I0(\processor/decode/instruction_reg_n_0_[6] ),
        .I1(\processor/id_shamt [3]),
        .I2(\processor/decode/instruction_reg_n_0_[5] ),
        .I3(\processor/id_rd_address [3]),
        .I4(\processor/decode/instruction_reg_n_0_[4] ),
        .I5(\processor/decode/instruction_reg_n_0_[3] ),
        .O(\immediate[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4000FFFF40000000)) 
    \immediate[4]_i_1 
       (.I0(\processor/decode/instruction_reg_n_0_[4] ),
        .I1(\processor/decode/instruction_reg_n_0_[6] ),
        .I2(\processor/id_shamt [4]),
        .I3(\processor/decode/instruction_reg_n_0_[5] ),
        .I4(\processor/decode/instruction_reg_n_0_ ),
        .I5(\immediate[4]_i_2_n_0 ),
        .O(\processor/id_immediate [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000008484F404)) 
    \immediate[4]_i_2 
       (.I0(\processor/decode/instruction_reg_n_0_[6] ),
        .I1(\processor/id_shamt [4]),
        .I2(\processor/decode/instruction_reg_n_0_[5] ),
        .I3(\processor/id_rd_address [4]),
        .I4(\processor/decode/instruction_reg_n_0_[4] ),
        .I5(\processor/decode/instruction_reg_n_0_[3] ),
        .O(\immediate[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \immediate_reg[0]_i_1 
       (.I0(immediate),
        .I1(\immediate[0]_i_3_n_0 ),
        .O(\processor/id_immediate [0]),
        .S(\processor/decode/instruction_reg_n_0_ ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \immediate_reg[11]_i_1 
       (.I0(\immediate[11]_i_2_n_0 ),
        .I1(\immediate[11]_i_3_n_0 ),
        .O(\processor/id_immediate [11]),
        .S(\processor/decode/instruction_reg_n_0_ ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \immediate_reg[12]_i_1 
       (.I0(\immediate[12]_i_2_n_0 ),
        .I1(\immediate[12]_i_3_n_0 ),
        .O(\processor/id_immediate [12]),
        .S(\processor/decode/instruction_reg_n_0_[3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \immediate_reg[13]_i_1 
       (.I0(\immediate[13]_i_2_n_0 ),
        .I1(\immediate[13]_i_3_n_0 ),
        .O(\processor/id_immediate [13]),
        .S(\processor/decode/instruction_reg_n_0_[3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \immediate_reg[14]_i_1 
       (.I0(\immediate[14]_i_2_n_0 ),
        .I1(\immediate[14]_i_3_n_0 ),
        .O(\processor/id_immediate [14]),
        .S(\processor/decode/instruction_reg_n_0_[3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \immediate_reg[15]_i_1 
       (.I0(\immediate[15]_i_2_n_0 ),
        .I1(\immediate[15]_i_3_n_0 ),
        .O(\processor/id_immediate [15]),
        .S(\processor/decode/instruction_reg_n_0_[3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \immediate_reg[16]_i_1 
       (.I0(\immediate[16]_i_2_n_0 ),
        .I1(\immediate[16]_i_3_n_0 ),
        .O(\processor/id_immediate [16]),
        .S(\processor/decode/instruction_reg_n_0_[3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \immediate_reg[17]_i_1 
       (.I0(\immediate[17]_i_2_n_0 ),
        .I1(\immediate[17]_i_3_n_0 ),
        .O(\processor/id_immediate [17]),
        .S(\processor/decode/instruction_reg_n_0_[3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \immediate_reg[18]_i_1 
       (.I0(\immediate[18]_i_2_n_0 ),
        .I1(\immediate[18]_i_3_n_0 ),
        .O(\processor/id_immediate [18]),
        .S(\processor/decode/instruction_reg_n_0_[3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \immediate_reg[19]_i_1 
       (.I0(\immediate[19]_i_2_n_0 ),
        .I1(\immediate[19]_i_3_n_0 ),
        .O(\processor/id_immediate [19]),
        .S(\processor/decode/instruction_reg_n_0_[3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \input_address_word[0]_i_1 
       (.I0(pc[2]),
        .I1(pc_next[2]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \input_address_word[1]_i_1 
       (.I0(pc[3]),
        .I1(pc_next[3]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB847000000000000)) 
    input_carry__0_i_1
       (.I0(\icache/tag_memory_reg_64_127_18_20_n_0 ),
        .I1(imem_address[10]),
        .I2(\icache/tag_memory_reg_0_63_18_20_n_0 ),
        .I3(imem_address[29]),
        .I4(input_carry__0_i_4_n_0),
        .I5(input_carry__0_i_5_n_0),
        .O(input_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB847000000000000)) 
    input_carry__0_i_2
       (.I0(\icache/tag_memory_reg_64_127_15_17_n_0 ),
        .I1(imem_address[10]),
        .I2(\icache/tag_memory_reg_0_63_15_17_n_0 ),
        .I3(imem_address[26]),
        .I4(input_carry__0_i_6_n_0),
        .I5(input_carry__0_i_7_n_0),
        .O(input_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB847000000000000)) 
    input_carry__0_i_3
       (.I0(\icache/tag_memory_reg_64_127_12_14_n_0 ),
        .I1(imem_address[10]),
        .I2(\icache/tag_memory_reg_0_63_12_14_n_0 ),
        .I3(imem_address[23]),
        .I4(input_carry__0_i_8_n_0),
        .I5(input_carry__0_i_9_n_0),
        .O(input_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hACACAC535353AC53)) 
    input_carry__0_i_4
       (.I0(pc[31]),
        .I1(pc_next[31]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/tag_memory_reg_0_63_18_20_n_2 ),
        .I4(imem_address[10]),
        .I5(\icache/tag_memory_reg_64_127_18_20_n_2 ),
        .O(input_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hACACAC535353AC53)) 
    input_carry__0_i_5
       (.I0(pc[30]),
        .I1(pc_next[30]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/tag_memory_reg_0_63_18_20_n_1 ),
        .I4(imem_address[10]),
        .I5(\icache/tag_memory_reg_64_127_18_20_n_1 ),
        .O(input_carry__0_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hACACAC535353AC53)) 
    input_carry__0_i_6
       (.I0(pc[28]),
        .I1(pc_next[28]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/tag_memory_reg_0_63_15_17_n_2 ),
        .I4(imem_address[10]),
        .I5(\icache/tag_memory_reg_64_127_15_17_n_2 ),
        .O(input_carry__0_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hACACAC535353AC53)) 
    input_carry__0_i_7
       (.I0(pc[27]),
        .I1(pc_next[27]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/tag_memory_reg_0_63_15_17_n_1 ),
        .I4(imem_address[10]),
        .I5(\icache/tag_memory_reg_64_127_15_17_n_1 ),
        .O(input_carry__0_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hACACAC535353AC53)) 
    input_carry__0_i_8
       (.I0(pc[25]),
        .I1(pc_next[25]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/tag_memory_reg_0_63_12_14_n_2 ),
        .I4(imem_address[10]),
        .I5(\icache/tag_memory_reg_64_127_12_14_n_2 ),
        .O(input_carry__0_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hACACAC535353AC53)) 
    input_carry__0_i_9
       (.I0(pc[24]),
        .I1(pc_next[24]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/tag_memory_reg_0_63_12_14_n_1 ),
        .I4(imem_address[10]),
        .I5(\icache/tag_memory_reg_64_127_12_14_n_1 ),
        .O(input_carry__0_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB847000000000000)) 
    input_carry_i_1
       (.I0(\icache/tag_memory_reg_64_127_9_11_n_0 ),
        .I1(imem_address[10]),
        .I2(\icache/tag_memory_reg_0_63_9_11_n_0 ),
        .I3(imem_address[20]),
        .I4(input_carry_i_5_n_0),
        .I5(input_carry_i_6_n_0),
        .O(input_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hACACAC535353AC53)) 
    input_carry_i_10
       (.I0(pc[15]),
        .I1(pc_next[15]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/tag_memory_reg_0_63_3_5_n_1 ),
        .I4(imem_address[10]),
        .I5(\icache/tag_memory_reg_64_127_3_5_n_1 ),
        .O(input_carry_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hACACAC535353AC53)) 
    input_carry_i_11
       (.I0(pc[13]),
        .I1(pc_next[13]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/tag_memory_reg_0_63_0_2_n_2 ),
        .I4(imem_address[10]),
        .I5(\icache/tag_memory_reg_64_127_0_2_n_2 ),
        .O(input_carry_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hACACAC535353AC53)) 
    input_carry_i_12
       (.I0(pc[12]),
        .I1(pc_next[12]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/tag_memory_reg_0_63_0_2_n_1 ),
        .I4(imem_address[10]),
        .I5(\icache/tag_memory_reg_64_127_0_2_n_1 ),
        .O(input_carry_i_12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB847000000000000)) 
    input_carry_i_2
       (.I0(\icache/tag_memory_reg_64_127_6_8_n_0 ),
        .I1(imem_address[10]),
        .I2(\icache/tag_memory_reg_0_63_6_8_n_0 ),
        .I3(imem_address[17]),
        .I4(input_carry_i_7_n_0),
        .I5(input_carry_i_8_n_0),
        .O(input_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB847000000000000)) 
    input_carry_i_3
       (.I0(\icache/tag_memory_reg_64_127_3_5_n_0 ),
        .I1(imem_address[10]),
        .I2(\icache/tag_memory_reg_0_63_3_5_n_0 ),
        .I3(imem_address[14]),
        .I4(input_carry_i_9_n_0),
        .I5(input_carry_i_10_n_0),
        .O(input_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB847000000000000)) 
    input_carry_i_4
       (.I0(\icache/tag_memory_reg_64_127_0_2_n_0 ),
        .I1(imem_address[10]),
        .I2(\icache/tag_memory_reg_0_63_0_2_n_0 ),
        .I3(imem_address[11]),
        .I4(input_carry_i_11_n_0),
        .I5(input_carry_i_12_n_0),
        .O(input_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hACACAC535353AC53)) 
    input_carry_i_5
       (.I0(pc[22]),
        .I1(pc_next[22]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/tag_memory_reg_0_63_9_11_n_2 ),
        .I4(imem_address[10]),
        .I5(\icache/tag_memory_reg_64_127_9_11_n_2 ),
        .O(input_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hACACAC535353AC53)) 
    input_carry_i_6
       (.I0(pc[21]),
        .I1(pc_next[21]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/tag_memory_reg_0_63_9_11_n_1 ),
        .I4(imem_address[10]),
        .I5(\icache/tag_memory_reg_64_127_9_11_n_1 ),
        .O(input_carry_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hACACAC535353AC53)) 
    input_carry_i_7
       (.I0(pc[19]),
        .I1(pc_next[19]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/tag_memory_reg_0_63_6_8_n_2 ),
        .I4(imem_address[10]),
        .I5(\icache/tag_memory_reg_64_127_6_8_n_2 ),
        .O(input_carry_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hACACAC535353AC53)) 
    input_carry_i_8
       (.I0(pc[18]),
        .I1(pc_next[18]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/tag_memory_reg_0_63_6_8_n_1 ),
        .I4(imem_address[10]),
        .I5(\icache/tag_memory_reg_64_127_6_8_n_1 ),
        .O(input_carry_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hACACAC535353AC53)) 
    input_carry_i_9
       (.I0(pc[16]),
        .I1(pc_next[16]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/tag_memory_reg_0_63_3_5_n_2 ),
        .I4(imem_address[10]),
        .I5(\icache/tag_memory_reg_64_127_3_5_n_2 ),
        .O(input_carry_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEEEEAEEEEEEEE)) 
    \instruction[31]_i_1 
       (.I0(reset),
        .I1(\processor/execute/exception_taken0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\mem_op[2]_i_5_n_0 ),
        .I4(\processor/fetch/cancel_fetch ),
        .I5(imem_ack),
        .O(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFE0002)) 
    \instruction[31]_i_3 
       (.I0(\icache/cache_hit ),
        .I1(\icache/state_reg_n_0_[2] ),
        .I2(\icache/state_reg_n_0_[1] ),
        .I3(\icache/state_reg_n_0_ ),
        .I4(\icache/read_ack ),
        .O(imem_ack));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[100]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[4]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(load_buffer));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[101]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[5]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[101]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[102]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[6]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[102]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[103]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[7]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[103]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[104]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[8]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[104]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[105]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[9]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[105]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[106]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[10]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[106]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[107]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[11]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[107]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[108]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[12]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[108]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[109]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[13]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[109]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[110]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[14]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[110]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[111]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[15]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[111]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[112]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[16]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[112]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[113]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[17]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[113]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[114]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[18]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[114]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[115]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[19]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[115]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[116]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[20]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[116]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[117]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[21]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[117]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[118]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[22]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[118]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[119]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[23]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[119]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[120]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[24]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[120]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[121]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[25]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[121]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[122]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[26]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[122]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[123]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[27]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[123]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[124]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[28]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[124]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[125]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[29]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[125]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[126]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[30]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[126]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0800000000000000)) 
    \load_buffer[127]_i_1 
       (.I0(\load_buffer[127]_i_3_n_0 ),
        .I1(\icache/cl_current_word_reg_n_0_[1] ),
        .I2(\icache/cl_current_word_reg_n_0_[2] ),
        .I3(\icache/cl_current_word_reg_n_0_ ),
        .I4(\icache/state_reg_n_0_ ),
        .I5(\icache/state_reg_n_0_[2] ),
        .O(\load_buffer[127]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[127]_i_2 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[31]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[127]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0008)) 
    \load_buffer[127]_i_3 
       (.I0(wb_ack_in),
        .I1(\arbiter/state [0]),
        .I2(\arbiter/state [1]),
        .I3(reset),
        .O(\load_buffer[127]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \load_buffer[31]_i_1 
       (.I0(\load_buffer[127]_i_3_n_0 ),
        .I1(\icache/cl_current_word_reg_n_0_ ),
        .I2(\icache/cl_current_word_reg_n_0_[2] ),
        .I3(\icache/cl_current_word_reg_n_0_[1] ),
        .I4(\icache/state_reg_n_0_ ),
        .I5(\icache/state_reg_n_0_[2] ),
        .O(\load_buffer[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \load_buffer[63]_i_1 
       (.I0(\load_buffer[127]_i_3_n_0 ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(\icache/cl_current_word_reg_n_0_ ),
        .I3(\icache/cl_current_word_reg_n_0_[1] ),
        .I4(\icache/state_reg_n_0_ ),
        .I5(\icache/state_reg_n_0_[2] ),
        .O(\load_buffer[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[64]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[0]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[64]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[65]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[1]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[65]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[66]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[2]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[66]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[67]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[3]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[67]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[68]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[4]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[68]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[69]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[5]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[69]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[70]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[6]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[70]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[71]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[7]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[71]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[72]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[8]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[72]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[73]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[9]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[73]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[74]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[10]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[74]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[75]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[11]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[75]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[76]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[12]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[76]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[77]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[13]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[77]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[78]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[14]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[78]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[79]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[15]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[79]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[80]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[16]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[80]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[81]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[17]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[81]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[82]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[18]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[82]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[83]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[19]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[83]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[84]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[20]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[84]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[85]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[21]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[85]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[86]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[22]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[86]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[87]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[23]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[87]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[88]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[24]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[88]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[89]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[25]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[89]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[90]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[26]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[90]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[91]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[27]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[91]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[92]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[28]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[92]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[93]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[29]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[93]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[94]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[30]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[94]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0008000000000000)) 
    \load_buffer[95]_i_1 
       (.I0(\load_buffer[127]_i_3_n_0 ),
        .I1(\icache/cl_current_word_reg_n_0_[1] ),
        .I2(\icache/cl_current_word_reg_n_0_ ),
        .I3(\icache/cl_current_word_reg_n_0_[2] ),
        .I4(\icache/state_reg_n_0_ ),
        .I5(\icache/state_reg_n_0_[2] ),
        .O(\load_buffer[95]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \load_buffer[95]_i_2 
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(wb_dat_in[31]),
        .I2(\arbiter/state [0]),
        .I3(\arbiter/state [1]),
        .I4(\icache/cl_current_word_reg_n_0_ ),
        .O(\load_buffer[95]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[96]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[0]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[96]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[97]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[1]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[97]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[98]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[2]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[98]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \load_buffer[99]_i_1 
       (.I0(\icache/cl_current_word_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(wb_dat_in[3]),
        .I3(\arbiter/state [0]),
        .I4(\arbiter/state [1]),
        .O(\load_buffer[99]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \mbadaddr[31]_i_1 
       (.I0(\processor/wb_exception ),
        .I1(reset),
        .O(\mbadaddr[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010000)) 
    \mem_op[0]_i_1 
       (.I0(\processor/decode/instruction_reg_n_0_ ),
        .I1(\processor/decode/instruction_reg_n_0_[6] ),
        .I2(\processor/decode/instruction_reg_n_0_[4] ),
        .I3(\processor/decode/instruction_reg_n_0_[3] ),
        .I4(mem_op),
        .O(\processor/id_mem_op [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFC8C)) 
    \mem_op[0]_i_2 
       (.I0(\processor/decode/instruction_reg_n_0_[5] ),
        .I1(\processor/id_csr_use_immediate ),
        .I2(\processor/id_funct3 [1]),
        .I3(\processor/id_funct3 [0]),
        .O(mem_op));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000010101)) 
    \mem_op[1]_i_1 
       (.I0(\processor/decode/instruction_reg_n_0_[6] ),
        .I1(\processor/decode/instruction_reg_n_0_[5] ),
        .I2(\processor/decode/instruction_reg_n_0_ ),
        .I3(\processor/id_funct3 [1]),
        .I4(\processor/id_funct3 [0]),
        .I5(\mem_op[1]_i_2_n_0 ),
        .O(\mem_op[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \mem_op[1]_i_2 
       (.I0(\processor/decode/instruction_reg_n_0_[4] ),
        .I1(\processor/decode/instruction_reg_n_0_[3] ),
        .O(\mem_op[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFE0)) 
    \mem_op[2]_i_1 
       (.I0(\mem_op[2]_i_4_n_0 ),
        .I1(\mem_op[2]_i_5_n_0 ),
        .I2(\processor/execute/exception_taken0 ),
        .I3(reset),
        .O(\processor/execute/rd_write_out0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_100 
       (.I0(\processor/ex_dmem_data_out [16]),
        .I1(\processor/execute/rs1_forwarded [16]),
        .I2(\processor/execute/rs1_forwarded [17]),
        .I3(\processor/ex_dmem_data_out [17]),
        .O(\mem_op[2]_i_100_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_101 
       (.I0(\processor/ex_dmem_data_out [22]),
        .I1(\processor/execute/rs1_forwarded [22]),
        .I2(\processor/ex_dmem_data_out [23]),
        .I3(\processor/execute/rs1_forwarded [23]),
        .O(\mem_op[2]_i_101_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_102 
       (.I0(\processor/ex_dmem_data_out [20]),
        .I1(\processor/execute/rs1_forwarded [20]),
        .I2(\processor/ex_dmem_data_out [21]),
        .I3(\processor/execute/rs1_forwarded [21]),
        .O(\mem_op[2]_i_102_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_103 
       (.I0(\processor/ex_dmem_data_out [18]),
        .I1(\processor/execute/rs1_forwarded [18]),
        .I2(\processor/ex_dmem_data_out [19]),
        .I3(\processor/execute/rs1_forwarded [19]),
        .O(\mem_op[2]_i_103_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_104 
       (.I0(\processor/ex_dmem_data_out [16]),
        .I1(\processor/execute/rs1_forwarded [16]),
        .I2(\processor/ex_dmem_data_out [17]),
        .I3(\processor/execute/rs1_forwarded [17]),
        .O(\mem_op[2]_i_104_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \mem_op[2]_i_105 
       (.I0(\processor/execute/rs1_forwarded [10]),
        .I1(\processor/ex_dmem_data_out [10]),
        .I2(\processor/execute/rs1_forwarded [11]),
        .I3(\processor/ex_dmem_data_out [11]),
        .I4(\processor/execute/rs1_forwarded [9]),
        .I5(\processor/ex_dmem_data_out [9]),
        .O(\mem_op[2]_i_105_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \mem_op[2]_i_106 
       (.I0(\processor/execute/rs1_forwarded [6]),
        .I1(\processor/ex_dmem_data_out [6]),
        .I2(\processor/ex_dmem_data_out [8]),
        .I3(\processor/execute/rs1_forwarded [8]),
        .I4(\processor/ex_dmem_data_out [7]),
        .I5(\processor/execute/rs1_forwarded [7]),
        .O(\mem_op[2]_i_106_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \mem_op[2]_i_107 
       (.I0(\processor/execute/rs1_forwarded [4]),
        .I1(\processor/ex_dmem_data_out [4]),
        .I2(\processor/execute/rs1_forwarded [5]),
        .I3(\processor/ex_dmem_data_out [5]),
        .I4(\processor/execute/rs1_forwarded [3]),
        .I5(\processor/ex_dmem_data_out [3]),
        .O(\mem_op[2]_i_107_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \mem_op[2]_i_108 
       (.I0(\processor/execute/rs1_forwarded [0]),
        .I1(\processor/ex_dmem_data_out [0]),
        .I2(\processor/ex_dmem_data_out [2]),
        .I3(\processor/execute/rs1_forwarded [2]),
        .I4(\processor/ex_dmem_data_out [1]),
        .I5(\processor/execute/rs1_forwarded [1]),
        .O(\mem_op[2]_i_108_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \mem_op[2]_i_109 
       (.I0(\processor/execute/rs1_forwarded [10]),
        .I1(\processor/ex_dmem_data_out [10]),
        .I2(\processor/execute/rs1_forwarded [11]),
        .I3(\processor/ex_dmem_data_out [11]),
        .I4(\processor/execute/rs1_forwarded [9]),
        .I5(\processor/ex_dmem_data_out [9]),
        .O(\mem_op[2]_i_109_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \mem_op[2]_i_110 
       (.I0(\processor/execute/rs1_forwarded [6]),
        .I1(\processor/ex_dmem_data_out [6]),
        .I2(\processor/ex_dmem_data_out [8]),
        .I3(\processor/execute/rs1_forwarded [8]),
        .I4(\processor/ex_dmem_data_out [7]),
        .I5(\processor/execute/rs1_forwarded [7]),
        .O(\mem_op[2]_i_110_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \mem_op[2]_i_111 
       (.I0(\processor/execute/rs1_forwarded [4]),
        .I1(\processor/ex_dmem_data_out [4]),
        .I2(\processor/execute/rs1_forwarded [5]),
        .I3(\processor/ex_dmem_data_out [5]),
        .I4(\processor/execute/rs1_forwarded [3]),
        .I5(\processor/ex_dmem_data_out [3]),
        .O(\mem_op[2]_i_111_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \mem_op[2]_i_112 
       (.I0(\processor/execute/rs1_forwarded [0]),
        .I1(\processor/ex_dmem_data_out [0]),
        .I2(\processor/ex_dmem_data_out [2]),
        .I3(\processor/execute/rs1_forwarded [2]),
        .I4(\processor/ex_dmem_data_out [1]),
        .I5(\processor/execute/rs1_forwarded [1]),
        .O(\mem_op[2]_i_112_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_114 
       (.I0(\processor/execute/rs1_forwarded [14]),
        .I1(\processor/ex_dmem_data_out [14]),
        .I2(\processor/ex_dmem_data_out [15]),
        .I3(\processor/execute/rs1_forwarded [15]),
        .O(\mem_op[2]_i_114_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_115 
       (.I0(\processor/execute/rs1_forwarded [12]),
        .I1(\processor/ex_dmem_data_out [12]),
        .I2(\processor/ex_dmem_data_out [13]),
        .I3(\processor/execute/rs1_forwarded [13]),
        .O(\mem_op[2]_i_115_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_116 
       (.I0(\processor/execute/rs1_forwarded [10]),
        .I1(\processor/ex_dmem_data_out [10]),
        .I2(\processor/ex_dmem_data_out [11]),
        .I3(\processor/execute/rs1_forwarded [11]),
        .O(\mem_op[2]_i_116_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_117 
       (.I0(\processor/execute/rs1_forwarded [8]),
        .I1(\processor/ex_dmem_data_out [8]),
        .I2(\processor/ex_dmem_data_out [9]),
        .I3(\processor/execute/rs1_forwarded [9]),
        .O(\mem_op[2]_i_117_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_118 
       (.I0(\processor/execute/rs1_forwarded [14]),
        .I1(\processor/ex_dmem_data_out [14]),
        .I2(\processor/execute/rs1_forwarded [15]),
        .I3(\processor/ex_dmem_data_out [15]),
        .O(\mem_op[2]_i_118_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_119 
       (.I0(\processor/execute/rs1_forwarded [12]),
        .I1(\processor/ex_dmem_data_out [12]),
        .I2(\processor/execute/rs1_forwarded [13]),
        .I3(\processor/ex_dmem_data_out [13]),
        .O(\mem_op[2]_i_119_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_120 
       (.I0(\processor/execute/rs1_forwarded [10]),
        .I1(\processor/ex_dmem_data_out [10]),
        .I2(\processor/execute/rs1_forwarded [11]),
        .I3(\processor/ex_dmem_data_out [11]),
        .O(\mem_op[2]_i_120_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_121 
       (.I0(\processor/execute/rs1_forwarded [8]),
        .I1(\processor/ex_dmem_data_out [8]),
        .I2(\processor/execute/rs1_forwarded [9]),
        .I3(\processor/ex_dmem_data_out [9]),
        .O(\mem_op[2]_i_121_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_123 
       (.I0(\processor/ex_dmem_data_out [14]),
        .I1(\processor/execute/rs1_forwarded [14]),
        .I2(\processor/execute/rs1_forwarded [15]),
        .I3(\processor/ex_dmem_data_out [15]),
        .O(\mem_op[2]_i_123_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_124 
       (.I0(\processor/ex_dmem_data_out [12]),
        .I1(\processor/execute/rs1_forwarded [12]),
        .I2(\processor/execute/rs1_forwarded [13]),
        .I3(\processor/ex_dmem_data_out [13]),
        .O(\mem_op[2]_i_124_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_125 
       (.I0(\processor/ex_dmem_data_out [10]),
        .I1(\processor/execute/rs1_forwarded [10]),
        .I2(\processor/execute/rs1_forwarded [11]),
        .I3(\processor/ex_dmem_data_out [11]),
        .O(\mem_op[2]_i_125_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_126 
       (.I0(\processor/ex_dmem_data_out [8]),
        .I1(\processor/execute/rs1_forwarded [8]),
        .I2(\processor/execute/rs1_forwarded [9]),
        .I3(\processor/ex_dmem_data_out [9]),
        .O(\mem_op[2]_i_126_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_127 
       (.I0(\processor/ex_dmem_data_out [14]),
        .I1(\processor/execute/rs1_forwarded [14]),
        .I2(\processor/ex_dmem_data_out [15]),
        .I3(\processor/execute/rs1_forwarded [15]),
        .O(\mem_op[2]_i_127_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_128 
       (.I0(\processor/ex_dmem_data_out [12]),
        .I1(\processor/execute/rs1_forwarded [12]),
        .I2(\processor/ex_dmem_data_out [13]),
        .I3(\processor/execute/rs1_forwarded [13]),
        .O(\mem_op[2]_i_128_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_129 
       (.I0(\processor/ex_dmem_data_out [10]),
        .I1(\processor/execute/rs1_forwarded [10]),
        .I2(\processor/ex_dmem_data_out [11]),
        .I3(\processor/execute/rs1_forwarded [11]),
        .O(\mem_op[2]_i_129_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_130 
       (.I0(\processor/ex_dmem_data_out [8]),
        .I1(\processor/execute/rs1_forwarded [8]),
        .I2(\processor/ex_dmem_data_out [9]),
        .I3(\processor/execute/rs1_forwarded [9]),
        .O(\mem_op[2]_i_130_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_132 
       (.I0(\processor/execute/rs1_forwarded [14]),
        .I1(\processor/ex_dmem_data_out [14]),
        .I2(\processor/ex_dmem_data_out [15]),
        .I3(\processor/execute/rs1_forwarded [15]),
        .O(\mem_op[2]_i_132_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_133 
       (.I0(\processor/execute/rs1_forwarded [12]),
        .I1(\processor/ex_dmem_data_out [12]),
        .I2(\processor/ex_dmem_data_out [13]),
        .I3(\processor/execute/rs1_forwarded [13]),
        .O(\mem_op[2]_i_133_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_134 
       (.I0(\processor/execute/rs1_forwarded [10]),
        .I1(\processor/ex_dmem_data_out [10]),
        .I2(\processor/ex_dmem_data_out [11]),
        .I3(\processor/execute/rs1_forwarded [11]),
        .O(\mem_op[2]_i_134_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_135 
       (.I0(\processor/execute/rs1_forwarded [8]),
        .I1(\processor/ex_dmem_data_out [8]),
        .I2(\processor/ex_dmem_data_out [9]),
        .I3(\processor/execute/rs1_forwarded [9]),
        .O(\mem_op[2]_i_135_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_136 
       (.I0(\processor/execute/rs1_forwarded [14]),
        .I1(\processor/ex_dmem_data_out [14]),
        .I2(\processor/execute/rs1_forwarded [15]),
        .I3(\processor/ex_dmem_data_out [15]),
        .O(\mem_op[2]_i_136_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_137 
       (.I0(\processor/execute/rs1_forwarded [12]),
        .I1(\processor/ex_dmem_data_out [12]),
        .I2(\processor/execute/rs1_forwarded [13]),
        .I3(\processor/ex_dmem_data_out [13]),
        .O(\mem_op[2]_i_137_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_138 
       (.I0(\processor/execute/rs1_forwarded [10]),
        .I1(\processor/ex_dmem_data_out [10]),
        .I2(\processor/execute/rs1_forwarded [11]),
        .I3(\processor/ex_dmem_data_out [11]),
        .O(\mem_op[2]_i_138_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_139 
       (.I0(\processor/execute/rs1_forwarded [8]),
        .I1(\processor/ex_dmem_data_out [8]),
        .I2(\processor/execute/rs1_forwarded [9]),
        .I3(\processor/ex_dmem_data_out [9]),
        .O(\mem_op[2]_i_139_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_141 
       (.I0(\processor/ex_dmem_data_out [14]),
        .I1(\processor/execute/rs1_forwarded [14]),
        .I2(\processor/execute/rs1_forwarded [15]),
        .I3(\processor/ex_dmem_data_out [15]),
        .O(\mem_op[2]_i_141_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_142 
       (.I0(\processor/ex_dmem_data_out [12]),
        .I1(\processor/execute/rs1_forwarded [12]),
        .I2(\processor/execute/rs1_forwarded [13]),
        .I3(\processor/ex_dmem_data_out [13]),
        .O(\mem_op[2]_i_142_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_143 
       (.I0(\processor/ex_dmem_data_out [10]),
        .I1(\processor/execute/rs1_forwarded [10]),
        .I2(\processor/execute/rs1_forwarded [11]),
        .I3(\processor/ex_dmem_data_out [11]),
        .O(\mem_op[2]_i_143_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_144 
       (.I0(\processor/ex_dmem_data_out [8]),
        .I1(\processor/execute/rs1_forwarded [8]),
        .I2(\processor/execute/rs1_forwarded [9]),
        .I3(\processor/ex_dmem_data_out [9]),
        .O(\mem_op[2]_i_144_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_145 
       (.I0(\processor/ex_dmem_data_out [14]),
        .I1(\processor/execute/rs1_forwarded [14]),
        .I2(\processor/ex_dmem_data_out [15]),
        .I3(\processor/execute/rs1_forwarded [15]),
        .O(\mem_op[2]_i_145_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_146 
       (.I0(\processor/ex_dmem_data_out [12]),
        .I1(\processor/execute/rs1_forwarded [12]),
        .I2(\processor/ex_dmem_data_out [13]),
        .I3(\processor/execute/rs1_forwarded [13]),
        .O(\mem_op[2]_i_146_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_147 
       (.I0(\processor/ex_dmem_data_out [10]),
        .I1(\processor/execute/rs1_forwarded [10]),
        .I2(\processor/ex_dmem_data_out [11]),
        .I3(\processor/execute/rs1_forwarded [11]),
        .O(\mem_op[2]_i_147_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_148 
       (.I0(\processor/ex_dmem_data_out [8]),
        .I1(\processor/execute/rs1_forwarded [8]),
        .I2(\processor/ex_dmem_data_out [9]),
        .I3(\processor/execute/rs1_forwarded [9]),
        .O(\mem_op[2]_i_148_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_149 
       (.I0(\processor/execute/rs1_forwarded [6]),
        .I1(\processor/ex_dmem_data_out [6]),
        .I2(\processor/ex_dmem_data_out [7]),
        .I3(\processor/execute/rs1_forwarded [7]),
        .O(\mem_op[2]_i_149_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_150 
       (.I0(\processor/execute/rs1_forwarded [4]),
        .I1(\processor/ex_dmem_data_out [4]),
        .I2(\processor/ex_dmem_data_out [5]),
        .I3(\processor/execute/rs1_forwarded [5]),
        .O(\mem_op[2]_i_150_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_151 
       (.I0(\processor/execute/rs1_forwarded [2]),
        .I1(\processor/ex_dmem_data_out [2]),
        .I2(\processor/ex_dmem_data_out [3]),
        .I3(\processor/execute/rs1_forwarded [3]),
        .O(\mem_op[2]_i_151_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_152 
       (.I0(\processor/execute/rs1_forwarded [0]),
        .I1(\processor/ex_dmem_data_out [0]),
        .I2(\processor/ex_dmem_data_out [1]),
        .I3(\processor/execute/rs1_forwarded [1]),
        .O(\mem_op[2]_i_152_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_153 
       (.I0(\processor/execute/rs1_forwarded [6]),
        .I1(\processor/ex_dmem_data_out [6]),
        .I2(\processor/execute/rs1_forwarded [7]),
        .I3(\processor/ex_dmem_data_out [7]),
        .O(\mem_op[2]_i_153_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_154 
       (.I0(\processor/execute/rs1_forwarded [4]),
        .I1(\processor/ex_dmem_data_out [4]),
        .I2(\processor/execute/rs1_forwarded [5]),
        .I3(\processor/ex_dmem_data_out [5]),
        .O(\mem_op[2]_i_154_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_155 
       (.I0(\processor/execute/rs1_forwarded [2]),
        .I1(\processor/ex_dmem_data_out [2]),
        .I2(\processor/execute/rs1_forwarded [3]),
        .I3(\processor/ex_dmem_data_out [3]),
        .O(\mem_op[2]_i_155_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_156 
       (.I0(\processor/execute/rs1_forwarded [0]),
        .I1(\processor/ex_dmem_data_out [0]),
        .I2(\processor/execute/rs1_forwarded [1]),
        .I3(\processor/ex_dmem_data_out [1]),
        .O(\mem_op[2]_i_156_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_157 
       (.I0(\processor/ex_dmem_data_out [6]),
        .I1(\processor/execute/rs1_forwarded [6]),
        .I2(\processor/execute/rs1_forwarded [7]),
        .I3(\processor/ex_dmem_data_out [7]),
        .O(\mem_op[2]_i_157_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_158 
       (.I0(\processor/ex_dmem_data_out [4]),
        .I1(\processor/execute/rs1_forwarded [4]),
        .I2(\processor/execute/rs1_forwarded [5]),
        .I3(\processor/ex_dmem_data_out [5]),
        .O(\mem_op[2]_i_158_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_159 
       (.I0(\processor/ex_dmem_data_out [2]),
        .I1(\processor/execute/rs1_forwarded [2]),
        .I2(\processor/execute/rs1_forwarded [3]),
        .I3(\processor/ex_dmem_data_out [3]),
        .O(\mem_op[2]_i_159_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_16 
       (.I0(\processor/ex_dmem_data_out [31]),
        .I1(\processor/execute/rs1_forwarded [31]),
        .I2(\processor/execute/rs1_forwarded [30]),
        .I3(\processor/ex_dmem_data_out [30]),
        .O(\mem_op[2]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_160 
       (.I0(\processor/ex_dmem_data_out [0]),
        .I1(\processor/execute/rs1_forwarded [0]),
        .I2(\processor/execute/rs1_forwarded [1]),
        .I3(\processor/ex_dmem_data_out [1]),
        .O(\mem_op[2]_i_160_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_161 
       (.I0(\processor/ex_dmem_data_out [6]),
        .I1(\processor/execute/rs1_forwarded [6]),
        .I2(\processor/ex_dmem_data_out [7]),
        .I3(\processor/execute/rs1_forwarded [7]),
        .O(\mem_op[2]_i_161_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_162 
       (.I0(\processor/ex_dmem_data_out [4]),
        .I1(\processor/execute/rs1_forwarded [4]),
        .I2(\processor/ex_dmem_data_out [5]),
        .I3(\processor/execute/rs1_forwarded [5]),
        .O(\mem_op[2]_i_162_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_163 
       (.I0(\processor/ex_dmem_data_out [2]),
        .I1(\processor/execute/rs1_forwarded [2]),
        .I2(\processor/ex_dmem_data_out [3]),
        .I3(\processor/execute/rs1_forwarded [3]),
        .O(\mem_op[2]_i_163_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_164 
       (.I0(\processor/ex_dmem_data_out [0]),
        .I1(\processor/execute/rs1_forwarded [0]),
        .I2(\processor/ex_dmem_data_out [1]),
        .I3(\processor/execute/rs1_forwarded [1]),
        .O(\mem_op[2]_i_164_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_165 
       (.I0(\processor/execute/rs1_forwarded [6]),
        .I1(\processor/ex_dmem_data_out [6]),
        .I2(\processor/ex_dmem_data_out [7]),
        .I3(\processor/execute/rs1_forwarded [7]),
        .O(\mem_op[2]_i_165_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_166 
       (.I0(\processor/execute/rs1_forwarded [4]),
        .I1(\processor/ex_dmem_data_out [4]),
        .I2(\processor/ex_dmem_data_out [5]),
        .I3(\processor/execute/rs1_forwarded [5]),
        .O(\mem_op[2]_i_166_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_167 
       (.I0(\processor/execute/rs1_forwarded [2]),
        .I1(\processor/ex_dmem_data_out [2]),
        .I2(\processor/ex_dmem_data_out [3]),
        .I3(\processor/execute/rs1_forwarded [3]),
        .O(\mem_op[2]_i_167_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_168 
       (.I0(\processor/execute/rs1_forwarded [0]),
        .I1(\processor/ex_dmem_data_out [0]),
        .I2(\processor/ex_dmem_data_out [1]),
        .I3(\processor/execute/rs1_forwarded [1]),
        .O(\mem_op[2]_i_168_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_169 
       (.I0(\processor/execute/rs1_forwarded [6]),
        .I1(\processor/ex_dmem_data_out [6]),
        .I2(\processor/execute/rs1_forwarded [7]),
        .I3(\processor/ex_dmem_data_out [7]),
        .O(\mem_op[2]_i_169_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \mem_op[2]_i_17 
       (.I0(\processor/execute/rs1_forwarded [28]),
        .I1(\processor/ex_dmem_data_out [28]),
        .I2(\processor/execute/rs1_forwarded [29]),
        .I3(\processor/ex_dmem_data_out [29]),
        .I4(\processor/execute/rs1_forwarded [27]),
        .I5(\processor/ex_dmem_data_out [27]),
        .O(\mem_op[2]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_170 
       (.I0(\processor/execute/rs1_forwarded [4]),
        .I1(\processor/ex_dmem_data_out [4]),
        .I2(\processor/execute/rs1_forwarded [5]),
        .I3(\processor/ex_dmem_data_out [5]),
        .O(\mem_op[2]_i_170_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_171 
       (.I0(\processor/execute/rs1_forwarded [2]),
        .I1(\processor/ex_dmem_data_out [2]),
        .I2(\processor/execute/rs1_forwarded [3]),
        .I3(\processor/ex_dmem_data_out [3]),
        .O(\mem_op[2]_i_171_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_172 
       (.I0(\processor/execute/rs1_forwarded [0]),
        .I1(\processor/ex_dmem_data_out [0]),
        .I2(\processor/execute/rs1_forwarded [1]),
        .I3(\processor/ex_dmem_data_out [1]),
        .O(\mem_op[2]_i_172_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_173 
       (.I0(\processor/ex_dmem_data_out [6]),
        .I1(\processor/execute/rs1_forwarded [6]),
        .I2(\processor/execute/rs1_forwarded [7]),
        .I3(\processor/ex_dmem_data_out [7]),
        .O(\mem_op[2]_i_173_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_174 
       (.I0(\processor/ex_dmem_data_out [4]),
        .I1(\processor/execute/rs1_forwarded [4]),
        .I2(\processor/execute/rs1_forwarded [5]),
        .I3(\processor/ex_dmem_data_out [5]),
        .O(\mem_op[2]_i_174_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_175 
       (.I0(\processor/ex_dmem_data_out [2]),
        .I1(\processor/execute/rs1_forwarded [2]),
        .I2(\processor/execute/rs1_forwarded [3]),
        .I3(\processor/ex_dmem_data_out [3]),
        .O(\mem_op[2]_i_175_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_176 
       (.I0(\processor/ex_dmem_data_out [0]),
        .I1(\processor/execute/rs1_forwarded [0]),
        .I2(\processor/execute/rs1_forwarded [1]),
        .I3(\processor/ex_dmem_data_out [1]),
        .O(\mem_op[2]_i_176_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_177 
       (.I0(\processor/ex_dmem_data_out [6]),
        .I1(\processor/execute/rs1_forwarded [6]),
        .I2(\processor/ex_dmem_data_out [7]),
        .I3(\processor/execute/rs1_forwarded [7]),
        .O(\mem_op[2]_i_177_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_178 
       (.I0(\processor/ex_dmem_data_out [4]),
        .I1(\processor/execute/rs1_forwarded [4]),
        .I2(\processor/ex_dmem_data_out [5]),
        .I3(\processor/execute/rs1_forwarded [5]),
        .O(\mem_op[2]_i_178_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_179 
       (.I0(\processor/ex_dmem_data_out [2]),
        .I1(\processor/execute/rs1_forwarded [2]),
        .I2(\processor/ex_dmem_data_out [3]),
        .I3(\processor/execute/rs1_forwarded [3]),
        .O(\mem_op[2]_i_179_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \mem_op[2]_i_18 
       (.I0(\processor/execute/rs1_forwarded [24]),
        .I1(\processor/ex_dmem_data_out [24]),
        .I2(\processor/ex_dmem_data_out [26]),
        .I3(\processor/execute/rs1_forwarded [26]),
        .I4(\processor/ex_dmem_data_out [25]),
        .I5(\processor/execute/rs1_forwarded [25]),
        .O(\mem_op[2]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_180 
       (.I0(\processor/ex_dmem_data_out [0]),
        .I1(\processor/execute/rs1_forwarded [0]),
        .I2(\processor/ex_dmem_data_out [1]),
        .I3(\processor/execute/rs1_forwarded [1]),
        .O(\mem_op[2]_i_180_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_20 
       (.I0(\processor/ex_dmem_data_out [31]),
        .I1(\processor/execute/rs1_forwarded [31]),
        .I2(\processor/execute/rs1_forwarded [30]),
        .I3(\processor/ex_dmem_data_out [30]),
        .O(\mem_op[2]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \mem_op[2]_i_21 
       (.I0(\processor/execute/rs1_forwarded [28]),
        .I1(\processor/ex_dmem_data_out [28]),
        .I2(\processor/execute/rs1_forwarded [29]),
        .I3(\processor/ex_dmem_data_out [29]),
        .I4(\processor/execute/rs1_forwarded [27]),
        .I5(\processor/ex_dmem_data_out [27]),
        .O(\mem_op[2]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \mem_op[2]_i_22 
       (.I0(\processor/execute/rs1_forwarded [24]),
        .I1(\processor/ex_dmem_data_out [24]),
        .I2(\processor/ex_dmem_data_out [26]),
        .I3(\processor/execute/rs1_forwarded [26]),
        .I4(\processor/ex_dmem_data_out [25]),
        .I5(\processor/execute/rs1_forwarded [25]),
        .O(\mem_op[2]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_24 
       (.I0(\processor/execute/rs1_forwarded [30]),
        .I1(\processor/ex_dmem_data_out [30]),
        .I2(\processor/ex_dmem_data_out [31]),
        .I3(\processor/execute/rs1_forwarded [31]),
        .O(\mem_op[2]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_25 
       (.I0(\processor/execute/rs1_forwarded [28]),
        .I1(\processor/ex_dmem_data_out [28]),
        .I2(\processor/ex_dmem_data_out [29]),
        .I3(\processor/execute/rs1_forwarded [29]),
        .O(\mem_op[2]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_26 
       (.I0(\processor/execute/rs1_forwarded [26]),
        .I1(\processor/ex_dmem_data_out [26]),
        .I2(\processor/ex_dmem_data_out [27]),
        .I3(\processor/execute/rs1_forwarded [27]),
        .O(\mem_op[2]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_27 
       (.I0(\processor/execute/rs1_forwarded [24]),
        .I1(\processor/ex_dmem_data_out [24]),
        .I2(\processor/ex_dmem_data_out [25]),
        .I3(\processor/execute/rs1_forwarded [25]),
        .O(\mem_op[2]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_28 
       (.I0(\processor/ex_dmem_data_out [31]),
        .I1(\processor/execute/rs1_forwarded [31]),
        .I2(\processor/execute/rs1_forwarded [30]),
        .I3(\processor/ex_dmem_data_out [30]),
        .O(\mem_op[2]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_29 
       (.I0(\processor/execute/rs1_forwarded [28]),
        .I1(\processor/ex_dmem_data_out [28]),
        .I2(\processor/execute/rs1_forwarded [29]),
        .I3(\processor/ex_dmem_data_out [29]),
        .O(\mem_op[2]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    \mem_op[2]_i_3 
       (.I0(\processor/decode/instruction_reg_n_0_[5] ),
        .I1(\processor/decode/instruction_reg_n_0_ ),
        .I2(\processor/id_csr_use_immediate ),
        .I3(\mem_op[2]_i_6_n_0 ),
        .O(\processor/id_mem_op [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_30 
       (.I0(\processor/execute/rs1_forwarded [26]),
        .I1(\processor/ex_dmem_data_out [26]),
        .I2(\processor/execute/rs1_forwarded [27]),
        .I3(\processor/ex_dmem_data_out [27]),
        .O(\mem_op[2]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_31 
       (.I0(\processor/execute/rs1_forwarded [24]),
        .I1(\processor/ex_dmem_data_out [24]),
        .I2(\processor/execute/rs1_forwarded [25]),
        .I3(\processor/ex_dmem_data_out [25]),
        .O(\mem_op[2]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_33 
       (.I0(\processor/ex_dmem_data_out [30]),
        .I1(\processor/execute/rs1_forwarded [30]),
        .I2(\processor/execute/rs1_forwarded [31]),
        .I3(\processor/ex_dmem_data_out [31]),
        .O(\mem_op[2]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_34 
       (.I0(\processor/ex_dmem_data_out [28]),
        .I1(\processor/execute/rs1_forwarded [28]),
        .I2(\processor/execute/rs1_forwarded [29]),
        .I3(\processor/ex_dmem_data_out [29]),
        .O(\mem_op[2]_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_35 
       (.I0(\processor/ex_dmem_data_out [26]),
        .I1(\processor/execute/rs1_forwarded [26]),
        .I2(\processor/execute/rs1_forwarded [27]),
        .I3(\processor/ex_dmem_data_out [27]),
        .O(\mem_op[2]_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_36 
       (.I0(\processor/ex_dmem_data_out [24]),
        .I1(\processor/execute/rs1_forwarded [24]),
        .I2(\processor/execute/rs1_forwarded [25]),
        .I3(\processor/ex_dmem_data_out [25]),
        .O(\mem_op[2]_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_37 
       (.I0(\processor/execute/rs1_forwarded [31]),
        .I1(\processor/ex_dmem_data_out [31]),
        .I2(\processor/ex_dmem_data_out [30]),
        .I3(\processor/execute/rs1_forwarded [30]),
        .O(\mem_op[2]_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_38 
       (.I0(\processor/ex_dmem_data_out [28]),
        .I1(\processor/execute/rs1_forwarded [28]),
        .I2(\processor/ex_dmem_data_out [29]),
        .I3(\processor/execute/rs1_forwarded [29]),
        .O(\mem_op[2]_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_39 
       (.I0(\processor/ex_dmem_data_out [26]),
        .I1(\processor/execute/rs1_forwarded [26]),
        .I2(\processor/ex_dmem_data_out [27]),
        .I3(\processor/execute/rs1_forwarded [27]),
        .O(\mem_op[2]_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h20222288)) 
    \mem_op[2]_i_4 
       (.I0(\processor/execute/exception_taken0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/execute/branch_condition ),
        .I3(\processor/ex_branch [1]),
        .I4(\processor/ex_branch [0]),
        .O(\mem_op[2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_40 
       (.I0(\processor/ex_dmem_data_out [24]),
        .I1(\processor/execute/rs1_forwarded [24]),
        .I2(\processor/ex_dmem_data_out [25]),
        .I3(\processor/execute/rs1_forwarded [25]),
        .O(\mem_op[2]_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_42 
       (.I0(\processor/execute/rs1_forwarded [30]),
        .I1(\processor/ex_dmem_data_out [30]),
        .I2(\processor/execute/rs1_forwarded [31]),
        .I3(\processor/ex_dmem_data_out [31]),
        .O(\mem_op[2]_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_43 
       (.I0(\processor/execute/rs1_forwarded [28]),
        .I1(\processor/ex_dmem_data_out [28]),
        .I2(\processor/ex_dmem_data_out [29]),
        .I3(\processor/execute/rs1_forwarded [29]),
        .O(\mem_op[2]_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_44 
       (.I0(\processor/execute/rs1_forwarded [26]),
        .I1(\processor/ex_dmem_data_out [26]),
        .I2(\processor/ex_dmem_data_out [27]),
        .I3(\processor/execute/rs1_forwarded [27]),
        .O(\mem_op[2]_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_45 
       (.I0(\processor/execute/rs1_forwarded [24]),
        .I1(\processor/ex_dmem_data_out [24]),
        .I2(\processor/ex_dmem_data_out [25]),
        .I3(\processor/execute/rs1_forwarded [25]),
        .O(\mem_op[2]_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_46 
       (.I0(\processor/execute/rs1_forwarded [31]),
        .I1(\processor/ex_dmem_data_out [31]),
        .I2(\processor/execute/rs1_forwarded [30]),
        .I3(\processor/ex_dmem_data_out [30]),
        .O(\mem_op[2]_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_47 
       (.I0(\processor/execute/rs1_forwarded [28]),
        .I1(\processor/ex_dmem_data_out [28]),
        .I2(\processor/execute/rs1_forwarded [29]),
        .I3(\processor/ex_dmem_data_out [29]),
        .O(\mem_op[2]_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_48 
       (.I0(\processor/execute/rs1_forwarded [26]),
        .I1(\processor/ex_dmem_data_out [26]),
        .I2(\processor/execute/rs1_forwarded [27]),
        .I3(\processor/ex_dmem_data_out [27]),
        .O(\mem_op[2]_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_49 
       (.I0(\processor/execute/rs1_forwarded [24]),
        .I1(\processor/ex_dmem_data_out [24]),
        .I2(\processor/execute/rs1_forwarded [25]),
        .I3(\processor/ex_dmem_data_out [25]),
        .O(\mem_op[2]_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAA8AAAA)) 
    \mem_op[2]_i_5 
       (.I0(\processor/execute/exception_taken0 ),
        .I1(\processor/execute/decode_exception ),
        .I2(\exception_context_out[cause][1]_i_2_n_0 ),
        .I3(\exception_context_out[cause][5]_i_2_n_0 ),
        .I4(\exception_context_out[cause][3]_i_3_n_0 ),
        .I5(\exception_context_out[cause][2]_i_2_n_0 ),
        .O(\mem_op[2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_51 
       (.I0(\processor/ex_dmem_data_out [30]),
        .I1(\processor/execute/rs1_forwarded [30]),
        .I2(\processor/ex_dmem_data_out [31]),
        .I3(\processor/execute/rs1_forwarded [31]),
        .O(\mem_op[2]_i_51_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_52 
       (.I0(\processor/ex_dmem_data_out [28]),
        .I1(\processor/execute/rs1_forwarded [28]),
        .I2(\processor/execute/rs1_forwarded [29]),
        .I3(\processor/ex_dmem_data_out [29]),
        .O(\mem_op[2]_i_52_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_53 
       (.I0(\processor/ex_dmem_data_out [26]),
        .I1(\processor/execute/rs1_forwarded [26]),
        .I2(\processor/execute/rs1_forwarded [27]),
        .I3(\processor/ex_dmem_data_out [27]),
        .O(\mem_op[2]_i_53_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_54 
       (.I0(\processor/ex_dmem_data_out [24]),
        .I1(\processor/execute/rs1_forwarded [24]),
        .I2(\processor/execute/rs1_forwarded [25]),
        .I3(\processor/ex_dmem_data_out [25]),
        .O(\mem_op[2]_i_54_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_55 
       (.I0(\processor/ex_dmem_data_out [31]),
        .I1(\processor/execute/rs1_forwarded [31]),
        .I2(\processor/ex_dmem_data_out [30]),
        .I3(\processor/execute/rs1_forwarded [30]),
        .O(\mem_op[2]_i_55_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_56 
       (.I0(\processor/ex_dmem_data_out [28]),
        .I1(\processor/execute/rs1_forwarded [28]),
        .I2(\processor/ex_dmem_data_out [29]),
        .I3(\processor/execute/rs1_forwarded [29]),
        .O(\mem_op[2]_i_56_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_57 
       (.I0(\processor/ex_dmem_data_out [26]),
        .I1(\processor/execute/rs1_forwarded [26]),
        .I2(\processor/ex_dmem_data_out [27]),
        .I3(\processor/execute/rs1_forwarded [27]),
        .O(\mem_op[2]_i_57_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_58 
       (.I0(\processor/ex_dmem_data_out [24]),
        .I1(\processor/execute/rs1_forwarded [24]),
        .I2(\processor/ex_dmem_data_out [25]),
        .I3(\processor/execute/rs1_forwarded [25]),
        .O(\mem_op[2]_i_58_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFEEE)) 
    \mem_op[2]_i_6 
       (.I0(\processor/decode/instruction_reg_n_0_[4] ),
        .I1(\processor/decode/instruction_reg_n_0_[6] ),
        .I2(\processor/id_funct3 [0]),
        .I3(\processor/id_funct3 [1]),
        .I4(\processor/decode/instruction_reg_n_0_[3] ),
        .O(\mem_op[2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \mem_op[2]_i_60 
       (.I0(\processor/execute/rs1_forwarded [22]),
        .I1(\processor/ex_dmem_data_out [22]),
        .I2(\processor/execute/rs1_forwarded [23]),
        .I3(\processor/ex_dmem_data_out [23]),
        .I4(\processor/execute/rs1_forwarded [21]),
        .I5(\processor/ex_dmem_data_out [21]),
        .O(\mem_op[2]_i_60_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \mem_op[2]_i_61 
       (.I0(\processor/execute/rs1_forwarded [18]),
        .I1(\processor/ex_dmem_data_out [18]),
        .I2(\processor/ex_dmem_data_out [20]),
        .I3(\processor/execute/rs1_forwarded [20]),
        .I4(\processor/ex_dmem_data_out [19]),
        .I5(\processor/execute/rs1_forwarded [19]),
        .O(\mem_op[2]_i_61_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \mem_op[2]_i_62 
       (.I0(\processor/execute/rs1_forwarded [16]),
        .I1(\processor/ex_dmem_data_out [16]),
        .I2(\processor/execute/rs1_forwarded [17]),
        .I3(\processor/ex_dmem_data_out [17]),
        .I4(\processor/execute/rs1_forwarded [15]),
        .I5(\processor/ex_dmem_data_out [15]),
        .O(\mem_op[2]_i_62_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \mem_op[2]_i_63 
       (.I0(\processor/execute/rs1_forwarded [12]),
        .I1(\processor/ex_dmem_data_out [12]),
        .I2(\processor/ex_dmem_data_out [14]),
        .I3(\processor/execute/rs1_forwarded [14]),
        .I4(\processor/ex_dmem_data_out [13]),
        .I5(\processor/execute/rs1_forwarded [13]),
        .O(\mem_op[2]_i_63_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \mem_op[2]_i_65 
       (.I0(\processor/execute/rs1_forwarded [22]),
        .I1(\processor/ex_dmem_data_out [22]),
        .I2(\processor/execute/rs1_forwarded [23]),
        .I3(\processor/ex_dmem_data_out [23]),
        .I4(\processor/execute/rs1_forwarded [21]),
        .I5(\processor/ex_dmem_data_out [21]),
        .O(\mem_op[2]_i_65_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \mem_op[2]_i_66 
       (.I0(\processor/execute/rs1_forwarded [18]),
        .I1(\processor/ex_dmem_data_out [18]),
        .I2(\processor/ex_dmem_data_out [20]),
        .I3(\processor/execute/rs1_forwarded [20]),
        .I4(\processor/ex_dmem_data_out [19]),
        .I5(\processor/execute/rs1_forwarded [19]),
        .O(\mem_op[2]_i_66_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \mem_op[2]_i_67 
       (.I0(\processor/execute/rs1_forwarded [16]),
        .I1(\processor/ex_dmem_data_out [16]),
        .I2(\processor/execute/rs1_forwarded [17]),
        .I3(\processor/ex_dmem_data_out [17]),
        .I4(\processor/execute/rs1_forwarded [15]),
        .I5(\processor/ex_dmem_data_out [15]),
        .O(\mem_op[2]_i_67_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \mem_op[2]_i_68 
       (.I0(\processor/execute/rs1_forwarded [12]),
        .I1(\processor/ex_dmem_data_out [12]),
        .I2(\processor/ex_dmem_data_out [14]),
        .I3(\processor/execute/rs1_forwarded [14]),
        .I4(\processor/ex_dmem_data_out [13]),
        .I5(\processor/execute/rs1_forwarded [13]),
        .O(\mem_op[2]_i_68_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA3A0A3A3A3A0A0A0)) 
    \mem_op[2]_i_7 
       (.I0(\mem_op[2]_i_8_n_0 ),
        .I1(\processor/execute/funct3 [1]),
        .I2(\processor/execute/funct3 [2]),
        .I3(\processor/execute/branch_comparator/data1 ),
        .I4(\processor/execute/funct3 [0]),
        .I5(\processor/execute/branch_comparator/data0 ),
        .O(\processor/execute/branch_condition ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_70 
       (.I0(\processor/execute/rs1_forwarded [22]),
        .I1(\processor/ex_dmem_data_out [22]),
        .I2(\processor/ex_dmem_data_out [23]),
        .I3(\processor/execute/rs1_forwarded [23]),
        .O(\mem_op[2]_i_70_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_71 
       (.I0(\processor/execute/rs1_forwarded [20]),
        .I1(\processor/ex_dmem_data_out [20]),
        .I2(\processor/ex_dmem_data_out [21]),
        .I3(\processor/execute/rs1_forwarded [21]),
        .O(\mem_op[2]_i_71_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_72 
       (.I0(\processor/execute/rs1_forwarded [18]),
        .I1(\processor/ex_dmem_data_out [18]),
        .I2(\processor/ex_dmem_data_out [19]),
        .I3(\processor/execute/rs1_forwarded [19]),
        .O(\mem_op[2]_i_72_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_73 
       (.I0(\processor/execute/rs1_forwarded [16]),
        .I1(\processor/ex_dmem_data_out [16]),
        .I2(\processor/ex_dmem_data_out [17]),
        .I3(\processor/execute/rs1_forwarded [17]),
        .O(\mem_op[2]_i_73_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_74 
       (.I0(\processor/execute/rs1_forwarded [22]),
        .I1(\processor/ex_dmem_data_out [22]),
        .I2(\processor/execute/rs1_forwarded [23]),
        .I3(\processor/ex_dmem_data_out [23]),
        .O(\mem_op[2]_i_74_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_75 
       (.I0(\processor/execute/rs1_forwarded [20]),
        .I1(\processor/ex_dmem_data_out [20]),
        .I2(\processor/execute/rs1_forwarded [21]),
        .I3(\processor/ex_dmem_data_out [21]),
        .O(\mem_op[2]_i_75_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_76 
       (.I0(\processor/execute/rs1_forwarded [18]),
        .I1(\processor/ex_dmem_data_out [18]),
        .I2(\processor/execute/rs1_forwarded [19]),
        .I3(\processor/ex_dmem_data_out [19]),
        .O(\mem_op[2]_i_76_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_77 
       (.I0(\processor/execute/rs1_forwarded [16]),
        .I1(\processor/ex_dmem_data_out [16]),
        .I2(\processor/execute/rs1_forwarded [17]),
        .I3(\processor/ex_dmem_data_out [17]),
        .O(\mem_op[2]_i_77_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_79 
       (.I0(\processor/ex_dmem_data_out [22]),
        .I1(\processor/execute/rs1_forwarded [22]),
        .I2(\processor/execute/rs1_forwarded [23]),
        .I3(\processor/ex_dmem_data_out [23]),
        .O(\mem_op[2]_i_79_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \mem_op[2]_i_8 
       (.I0(\processor/execute/branch_comparator/data5 ),
        .I1(\processor/execute/branch_comparator/data4 ),
        .I2(\processor/execute/funct3 [1]),
        .I3(\processor/execute/branch_comparator/data3 ),
        .I4(\processor/execute/funct3 [0]),
        .I5(\processor/execute/branch_comparator/data2 ),
        .O(\mem_op[2]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_80 
       (.I0(\processor/ex_dmem_data_out [20]),
        .I1(\processor/execute/rs1_forwarded [20]),
        .I2(\processor/execute/rs1_forwarded [21]),
        .I3(\processor/ex_dmem_data_out [21]),
        .O(\mem_op[2]_i_80_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_81 
       (.I0(\processor/ex_dmem_data_out [18]),
        .I1(\processor/execute/rs1_forwarded [18]),
        .I2(\processor/execute/rs1_forwarded [19]),
        .I3(\processor/ex_dmem_data_out [19]),
        .O(\mem_op[2]_i_81_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_82 
       (.I0(\processor/ex_dmem_data_out [16]),
        .I1(\processor/execute/rs1_forwarded [16]),
        .I2(\processor/execute/rs1_forwarded [17]),
        .I3(\processor/ex_dmem_data_out [17]),
        .O(\mem_op[2]_i_82_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_83 
       (.I0(\processor/ex_dmem_data_out [22]),
        .I1(\processor/execute/rs1_forwarded [22]),
        .I2(\processor/ex_dmem_data_out [23]),
        .I3(\processor/execute/rs1_forwarded [23]),
        .O(\mem_op[2]_i_83_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_84 
       (.I0(\processor/ex_dmem_data_out [20]),
        .I1(\processor/execute/rs1_forwarded [20]),
        .I2(\processor/ex_dmem_data_out [21]),
        .I3(\processor/execute/rs1_forwarded [21]),
        .O(\mem_op[2]_i_84_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_85 
       (.I0(\processor/ex_dmem_data_out [18]),
        .I1(\processor/execute/rs1_forwarded [18]),
        .I2(\processor/ex_dmem_data_out [19]),
        .I3(\processor/execute/rs1_forwarded [19]),
        .O(\mem_op[2]_i_85_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_86 
       (.I0(\processor/ex_dmem_data_out [16]),
        .I1(\processor/execute/rs1_forwarded [16]),
        .I2(\processor/ex_dmem_data_out [17]),
        .I3(\processor/execute/rs1_forwarded [17]),
        .O(\mem_op[2]_i_86_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_88 
       (.I0(\processor/execute/rs1_forwarded [22]),
        .I1(\processor/ex_dmem_data_out [22]),
        .I2(\processor/ex_dmem_data_out [23]),
        .I3(\processor/execute/rs1_forwarded [23]),
        .O(\mem_op[2]_i_88_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_89 
       (.I0(\processor/execute/rs1_forwarded [20]),
        .I1(\processor/ex_dmem_data_out [20]),
        .I2(\processor/ex_dmem_data_out [21]),
        .I3(\processor/execute/rs1_forwarded [21]),
        .O(\mem_op[2]_i_89_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_90 
       (.I0(\processor/execute/rs1_forwarded [18]),
        .I1(\processor/ex_dmem_data_out [18]),
        .I2(\processor/ex_dmem_data_out [19]),
        .I3(\processor/execute/rs1_forwarded [19]),
        .O(\mem_op[2]_i_90_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_91 
       (.I0(\processor/execute/rs1_forwarded [16]),
        .I1(\processor/ex_dmem_data_out [16]),
        .I2(\processor/ex_dmem_data_out [17]),
        .I3(\processor/execute/rs1_forwarded [17]),
        .O(\mem_op[2]_i_91_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_92 
       (.I0(\processor/execute/rs1_forwarded [22]),
        .I1(\processor/ex_dmem_data_out [22]),
        .I2(\processor/execute/rs1_forwarded [23]),
        .I3(\processor/ex_dmem_data_out [23]),
        .O(\mem_op[2]_i_92_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_93 
       (.I0(\processor/execute/rs1_forwarded [20]),
        .I1(\processor/ex_dmem_data_out [20]),
        .I2(\processor/execute/rs1_forwarded [21]),
        .I3(\processor/ex_dmem_data_out [21]),
        .O(\mem_op[2]_i_93_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_94 
       (.I0(\processor/execute/rs1_forwarded [18]),
        .I1(\processor/ex_dmem_data_out [18]),
        .I2(\processor/execute/rs1_forwarded [19]),
        .I3(\processor/ex_dmem_data_out [19]),
        .O(\mem_op[2]_i_94_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \mem_op[2]_i_95 
       (.I0(\processor/execute/rs1_forwarded [16]),
        .I1(\processor/ex_dmem_data_out [16]),
        .I2(\processor/execute/rs1_forwarded [17]),
        .I3(\processor/ex_dmem_data_out [17]),
        .O(\mem_op[2]_i_95_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_97 
       (.I0(\processor/ex_dmem_data_out [22]),
        .I1(\processor/execute/rs1_forwarded [22]),
        .I2(\processor/execute/rs1_forwarded [23]),
        .I3(\processor/ex_dmem_data_out [23]),
        .O(\mem_op[2]_i_97_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_98 
       (.I0(\processor/ex_dmem_data_out [20]),
        .I1(\processor/execute/rs1_forwarded [20]),
        .I2(\processor/execute/rs1_forwarded [21]),
        .I3(\processor/ex_dmem_data_out [21]),
        .O(\mem_op[2]_i_98_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \mem_op[2]_i_99 
       (.I0(\processor/ex_dmem_data_out [18]),
        .I1(\processor/execute/rs1_forwarded [18]),
        .I2(\processor/execute/rs1_forwarded [19]),
        .I3(\processor/ex_dmem_data_out [19]),
        .O(\mem_op[2]_i_99_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mem_op_reg[2]_i_10 
       (.CI(\mem_op_reg[2]_i_19_n_0 ),
        .CO({\mem_op_reg[2]_i_10_n_0 ,\processor/execute/branch_comparator/data0 ,\mem_op_reg[2]_i_10_n_2 ,\mem_op_reg[2]_i_10_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const0>__0__0 ,\mem_op[2]_i_20_n_0 ,\mem_op[2]_i_21_n_0 ,\mem_op[2]_i_22_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mem_op_reg[2]_i_11 
       (.CI(\mem_op_reg[2]_i_23_n_0 ),
        .CO({\processor/execute/branch_comparator/data5 ,\mem_op_reg[2]_i_11_n_1 ,\mem_op_reg[2]_i_11_n_2 ,\mem_op_reg[2]_i_11_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\mem_op[2]_i_24_n_0 ,\mem_op[2]_i_25_n_0 ,\mem_op[2]_i_26_n_0 ,\mem_op[2]_i_27_n_0 }),
        .S({\mem_op[2]_i_28_n_0 ,\mem_op[2]_i_29_n_0 ,\mem_op[2]_i_30_n_0 ,\mem_op[2]_i_31_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mem_op_reg[2]_i_113 
       (.CI(\<const0>__0__0 ),
        .CO(mem_op_reg),
        .CYINIT(\<const1>__0__0 ),
        .DI({\mem_op[2]_i_149_n_0 ,\mem_op[2]_i_150_n_0 ,\mem_op[2]_i_151_n_0 ,\mem_op[2]_i_152_n_0 }),
        .S({\mem_op[2]_i_153_n_0 ,\mem_op[2]_i_154_n_0 ,\mem_op[2]_i_155_n_0 ,\mem_op[2]_i_156_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mem_op_reg[2]_i_12 
       (.CI(\mem_op_reg[2]_i_32_n_0 ),
        .CO({\processor/execute/branch_comparator/data4 ,\mem_op_reg[2]_i_12_n_1 ,\mem_op_reg[2]_i_12_n_2 ,\mem_op_reg[2]_i_12_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\mem_op[2]_i_33_n_0 ,\mem_op[2]_i_34_n_0 ,\mem_op[2]_i_35_n_0 ,\mem_op[2]_i_36_n_0 }),
        .S({\mem_op[2]_i_37_n_0 ,\mem_op[2]_i_38_n_0 ,\mem_op[2]_i_39_n_0 ,\mem_op[2]_i_40_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mem_op_reg[2]_i_122 
       (.CI(\<const0>__0__0 ),
        .CO({\mem_op_reg[2]_i_122_n_0 ,\mem_op_reg[2]_i_122_n_1 ,\mem_op_reg[2]_i_122_n_2 ,\mem_op_reg[2]_i_122_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\mem_op[2]_i_157_n_0 ,\mem_op[2]_i_158_n_0 ,\mem_op[2]_i_159_n_0 ,\mem_op[2]_i_160_n_0 }),
        .S({\mem_op[2]_i_161_n_0 ,\mem_op[2]_i_162_n_0 ,\mem_op[2]_i_163_n_0 ,\mem_op[2]_i_164_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mem_op_reg[2]_i_13 
       (.CI(\mem_op_reg[2]_i_41_n_0 ),
        .CO({\processor/execute/branch_comparator/data3 ,\mem_op_reg[2]_i_13_n_1 ,\mem_op_reg[2]_i_13_n_2 ,\mem_op_reg[2]_i_13_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\mem_op[2]_i_42_n_0 ,\mem_op[2]_i_43_n_0 ,\mem_op[2]_i_44_n_0 ,\mem_op[2]_i_45_n_0 }),
        .S({\mem_op[2]_i_46_n_0 ,\mem_op[2]_i_47_n_0 ,\mem_op[2]_i_48_n_0 ,\mem_op[2]_i_49_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mem_op_reg[2]_i_131 
       (.CI(\<const0>__0__0 ),
        .CO({\mem_op_reg[2]_i_131_n_0 ,\mem_op_reg[2]_i_131_n_1 ,\mem_op_reg[2]_i_131_n_2 ,\mem_op_reg[2]_i_131_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\mem_op[2]_i_165_n_0 ,\mem_op[2]_i_166_n_0 ,\mem_op[2]_i_167_n_0 ,\mem_op[2]_i_168_n_0 }),
        .S({\mem_op[2]_i_169_n_0 ,\mem_op[2]_i_170_n_0 ,\mem_op[2]_i_171_n_0 ,\mem_op[2]_i_172_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mem_op_reg[2]_i_14 
       (.CI(\mem_op_reg[2]_i_50_n_0 ),
        .CO({\processor/execute/branch_comparator/data2 ,\mem_op_reg[2]_i_14_n_1 ,\mem_op_reg[2]_i_14_n_2 ,\mem_op_reg[2]_i_14_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\mem_op[2]_i_51_n_0 ,\mem_op[2]_i_52_n_0 ,\mem_op[2]_i_53_n_0 ,\mem_op[2]_i_54_n_0 }),
        .S({\mem_op[2]_i_55_n_0 ,\mem_op[2]_i_56_n_0 ,\mem_op[2]_i_57_n_0 ,\mem_op[2]_i_58_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mem_op_reg[2]_i_140 
       (.CI(\<const0>__0__0 ),
        .CO({\mem_op_reg[2]_i_140_n_0 ,\mem_op_reg[2]_i_140_n_1 ,\mem_op_reg[2]_i_140_n_2 ,\mem_op_reg[2]_i_140_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\mem_op[2]_i_173_n_0 ,\mem_op[2]_i_174_n_0 ,\mem_op[2]_i_175_n_0 ,\mem_op[2]_i_176_n_0 }),
        .S({\mem_op[2]_i_177_n_0 ,\mem_op[2]_i_178_n_0 ,\mem_op[2]_i_179_n_0 ,\mem_op[2]_i_180_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mem_op_reg[2]_i_15 
       (.CI(\mem_op_reg[2]_i_59_n_0 ),
        .CO({\mem_op_reg[2]_i_15_n_0 ,\mem_op_reg[2]_i_15_n_1 ,\mem_op_reg[2]_i_15_n_2 ,\mem_op_reg[2]_i_15_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\mem_op[2]_i_60_n_0 ,\mem_op[2]_i_61_n_0 ,\mem_op[2]_i_62_n_0 ,\mem_op[2]_i_63_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mem_op_reg[2]_i_19 
       (.CI(\mem_op_reg[2]_i_64_n_0 ),
        .CO({\mem_op_reg[2]_i_19_n_0 ,\mem_op_reg[2]_i_19_n_1 ,\mem_op_reg[2]_i_19_n_2 ,\mem_op_reg[2]_i_19_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\mem_op[2]_i_65_n_0 ,\mem_op[2]_i_66_n_0 ,\mem_op[2]_i_67_n_0 ,\mem_op[2]_i_68_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mem_op_reg[2]_i_23 
       (.CI(\mem_op_reg[2]_i_69_n_0 ),
        .CO({\mem_op_reg[2]_i_23_n_0 ,\mem_op_reg[2]_i_23_n_1 ,\mem_op_reg[2]_i_23_n_2 ,\mem_op_reg[2]_i_23_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\mem_op[2]_i_70_n_0 ,\mem_op[2]_i_71_n_0 ,\mem_op[2]_i_72_n_0 ,\mem_op[2]_i_73_n_0 }),
        .S({\mem_op[2]_i_74_n_0 ,\mem_op[2]_i_75_n_0 ,\mem_op[2]_i_76_n_0 ,\mem_op[2]_i_77_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mem_op_reg[2]_i_32 
       (.CI(\mem_op_reg[2]_i_78_n_0 ),
        .CO({\mem_op_reg[2]_i_32_n_0 ,\mem_op_reg[2]_i_32_n_1 ,\mem_op_reg[2]_i_32_n_2 ,\mem_op_reg[2]_i_32_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\mem_op[2]_i_79_n_0 ,\mem_op[2]_i_80_n_0 ,\mem_op[2]_i_81_n_0 ,\mem_op[2]_i_82_n_0 }),
        .S({\mem_op[2]_i_83_n_0 ,\mem_op[2]_i_84_n_0 ,\mem_op[2]_i_85_n_0 ,\mem_op[2]_i_86_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mem_op_reg[2]_i_41 
       (.CI(\mem_op_reg[2]_i_87_n_0 ),
        .CO({\mem_op_reg[2]_i_41_n_0 ,\mem_op_reg[2]_i_41_n_1 ,\mem_op_reg[2]_i_41_n_2 ,\mem_op_reg[2]_i_41_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\mem_op[2]_i_88_n_0 ,\mem_op[2]_i_89_n_0 ,\mem_op[2]_i_90_n_0 ,\mem_op[2]_i_91_n_0 }),
        .S({\mem_op[2]_i_92_n_0 ,\mem_op[2]_i_93_n_0 ,\mem_op[2]_i_94_n_0 ,\mem_op[2]_i_95_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mem_op_reg[2]_i_50 
       (.CI(\mem_op_reg[2]_i_96_n_0 ),
        .CO({\mem_op_reg[2]_i_50_n_0 ,\mem_op_reg[2]_i_50_n_1 ,\mem_op_reg[2]_i_50_n_2 ,\mem_op_reg[2]_i_50_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\mem_op[2]_i_97_n_0 ,\mem_op[2]_i_98_n_0 ,\mem_op[2]_i_99_n_0 ,\mem_op[2]_i_100_n_0 }),
        .S({\mem_op[2]_i_101_n_0 ,\mem_op[2]_i_102_n_0 ,\mem_op[2]_i_103_n_0 ,\mem_op[2]_i_104_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mem_op_reg[2]_i_59 
       (.CI(\<const0>__0__0 ),
        .CO({\mem_op_reg[2]_i_59_n_0 ,\mem_op_reg[2]_i_59_n_1 ,\mem_op_reg[2]_i_59_n_2 ,\mem_op_reg[2]_i_59_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\mem_op[2]_i_105_n_0 ,\mem_op[2]_i_106_n_0 ,\mem_op[2]_i_107_n_0 ,\mem_op[2]_i_108_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mem_op_reg[2]_i_64 
       (.CI(\<const0>__0__0 ),
        .CO({\mem_op_reg[2]_i_64_n_0 ,\mem_op_reg[2]_i_64_n_1 ,\mem_op_reg[2]_i_64_n_2 ,\mem_op_reg[2]_i_64_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\mem_op[2]_i_109_n_0 ,\mem_op[2]_i_110_n_0 ,\mem_op[2]_i_111_n_0 ,\mem_op[2]_i_112_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mem_op_reg[2]_i_69 
       (.CI(mem_op_reg[3]),
        .CO({\mem_op_reg[2]_i_69_n_0 ,\mem_op_reg[2]_i_69_n_1 ,\mem_op_reg[2]_i_69_n_2 ,\mem_op_reg[2]_i_69_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\mem_op[2]_i_114_n_0 ,\mem_op[2]_i_115_n_0 ,\mem_op[2]_i_116_n_0 ,\mem_op[2]_i_117_n_0 }),
        .S({\mem_op[2]_i_118_n_0 ,\mem_op[2]_i_119_n_0 ,\mem_op[2]_i_120_n_0 ,\mem_op[2]_i_121_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mem_op_reg[2]_i_78 
       (.CI(\mem_op_reg[2]_i_122_n_0 ),
        .CO({\mem_op_reg[2]_i_78_n_0 ,\mem_op_reg[2]_i_78_n_1 ,\mem_op_reg[2]_i_78_n_2 ,\mem_op_reg[2]_i_78_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\mem_op[2]_i_123_n_0 ,\mem_op[2]_i_124_n_0 ,\mem_op[2]_i_125_n_0 ,\mem_op[2]_i_126_n_0 }),
        .S({\mem_op[2]_i_127_n_0 ,\mem_op[2]_i_128_n_0 ,\mem_op[2]_i_129_n_0 ,\mem_op[2]_i_130_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mem_op_reg[2]_i_87 
       (.CI(\mem_op_reg[2]_i_131_n_0 ),
        .CO({\mem_op_reg[2]_i_87_n_0 ,\mem_op_reg[2]_i_87_n_1 ,\mem_op_reg[2]_i_87_n_2 ,\mem_op_reg[2]_i_87_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\mem_op[2]_i_132_n_0 ,\mem_op[2]_i_133_n_0 ,\mem_op[2]_i_134_n_0 ,\mem_op[2]_i_135_n_0 }),
        .S({\mem_op[2]_i_136_n_0 ,\mem_op[2]_i_137_n_0 ,\mem_op[2]_i_138_n_0 ,\mem_op[2]_i_139_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mem_op_reg[2]_i_9 
       (.CI(\mem_op_reg[2]_i_15_n_0 ),
        .CO({\mem_op_reg[2]_i_9_n_0 ,\processor/execute/branch_comparator/data1 ,\mem_op_reg[2]_i_9_n_2 ,\mem_op_reg[2]_i_9_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\<const0>__0__0 ,\mem_op[2]_i_16_n_0 ,\mem_op[2]_i_17_n_0 ,\mem_op[2]_i_18_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mem_op_reg[2]_i_96 
       (.CI(\mem_op_reg[2]_i_140_n_0 ),
        .CO({\mem_op_reg[2]_i_96_n_0 ,\mem_op_reg[2]_i_96_n_1 ,\mem_op_reg[2]_i_96_n_2 ,\mem_op_reg[2]_i_96_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\mem_op[2]_i_141_n_0 ,\mem_op[2]_i_142_n_0 ,\mem_op[2]_i_143_n_0 ,\mem_op[2]_i_144_n_0 }),
        .S({\mem_op[2]_i_145_n_0 ,\mem_op[2]_i_146_n_0 ,\mem_op[2]_i_147_n_0 ,\mem_op[2]_i_148_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \mem_size[0]_i_1 
       (.I0(\mem_size[0]_i_2_n_0 ),
        .I1(\processor/id_funct3 [0]),
        .I2(\processor/decode/instruction_reg_n_0_[3] ),
        .I3(\mem_size[0]_i_3_n_0 ),
        .I4(\processor/decode/instruction_reg_n_0_ ),
        .I5(\processor/decode/instruction_reg_n_0_[4] ),
        .O(\processor/id_mem_size ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \mem_size[0]_i_2 
       (.I0(\processor/decode/instruction_reg_n_0_[6] ),
        .I1(\processor/id_funct3 [1]),
        .O(\mem_size[0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \mem_size[0]_i_3 
       (.I0(\processor/decode/instruction_reg_n_0_[5] ),
        .I1(\processor/id_csr_use_immediate ),
        .O(\mem_size[0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    \mem_size[1]_i_1 
       (.I0(\mem_op[2]_i_4_n_0 ),
        .I1(\mem_op[2]_i_5_n_0 ),
        .I2(\processor/execute/exception_taken0 ),
        .I3(reset),
        .O(\mem_size[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEA)) 
    \mem_size[1]_i_2 
       (.I0(\processor/decode/instruction_reg_n_0_ ),
        .I1(\processor/id_csr_use_immediate ),
        .I2(\processor/decode/instruction_reg_n_0_[5] ),
        .I3(\mem_op[1]_i_2_n_0 ),
        .I4(\processor/id_funct3 [1]),
        .I5(\processor/decode/instruction_reg_n_0_[6] ),
        .O(\mem_size[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \mepc[31]_i_1 
       (.I0(\processor/csr_unit/tohost_data1__0 ),
        .I1(\mtime_compare[31]_i_3_n_0 ),
        .I2(\processor/wb_csr_address [5]),
        .I3(\processor/wb_csr_address [1]),
        .I4(\processor/wb_csr_address [0]),
        .I5(\mepc[31]_i_2_n_0 ),
        .O(\mepc[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFEFF)) 
    \mepc[31]_i_2 
       (.I0(\processor/wb_csr_address [3]),
        .I1(\processor/wb_csr_address [4]),
        .I2(\processor/wb_csr_address [2]),
        .I3(\processor/wb_csr_address [6]),
        .O(\mepc[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \mie[31]_i_1 
       (.I0(\processor/csr_unit/tohost_data1__0 ),
        .I1(\mtime_compare[31]_i_3_n_0 ),
        .I2(\processor/wb_csr_address [6]),
        .I3(\processor/wb_csr_address [5]),
        .I4(\processor/wb_csr_address [2]),
        .I5(\mie[31]_i_2_n_0 ),
        .O(mie));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \mie[31]_i_2 
       (.I0(\processor/wb_csr_address [1]),
        .I1(\processor/wb_csr_address [0]),
        .I2(\processor/wb_csr_address [3]),
        .I3(\processor/wb_csr_address [4]),
        .O(\mie[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000E00)) 
    \mscratch[31]_i_1 
       (.I0(\processor/wb_csr_write [0]),
        .I1(\processor/wb_csr_write [1]),
        .I2(reset),
        .I3(\processor/csr_unit/mscratch__4 ),
        .I4(\mtime_compare[31]_i_3_n_0 ),
        .O(\mscratch[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000001000000000)) 
    \mscratch[31]_i_2 
       (.I0(\processor/wb_csr_address [5]),
        .I1(\processor/wb_csr_address [0]),
        .I2(\processor/wb_csr_address [6]),
        .I3(\processor/wb_csr_address [2]),
        .I4(\processor/wb_csr_address [1]),
        .I5(\mtime_compare[31]_i_4_n_0 ),
        .O(\processor/csr_unit/mscratch__4 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000E00)) 
    \mtime_compare[31]_i_1 
       (.I0(\processor/wb_csr_write [0]),
        .I1(\processor/wb_csr_write [1]),
        .I2(reset),
        .I3(\processor/csr_unit/mtime_compare__4 ),
        .I4(\mtime_compare[31]_i_3_n_0 ),
        .O(\mtime_compare[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \mtime_compare[31]_i_2 
       (.I0(\processor/wb_csr_address [1]),
        .I1(\processor/wb_csr_address [6]),
        .I2(\processor/wb_csr_address [0]),
        .I3(\processor/wb_csr_address [5]),
        .I4(\processor/wb_csr_address [2]),
        .I5(\mtime_compare[31]_i_4_n_0 ),
        .O(\processor/csr_unit/mtime_compare__4 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFDFFFF)) 
    \mtime_compare[31]_i_3 
       (.I0(\processor/wb_csr_address [9]),
        .I1(\processor/wb_csr_address [11]),
        .I2(\processor/wb_csr_address [10]),
        .I3(\processor/wb_csr_address [7]),
        .I4(\processor/wb_csr_address [8]),
        .O(\mtime_compare[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \mtime_compare[31]_i_4 
       (.I0(\processor/wb_csr_address [4]),
        .I1(\processor/wb_csr_address [3]),
        .O(\mtime_compare[31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \mtvec[31]_i_1 
       (.I0(\processor/csr_unit/tohost_data1__0 ),
        .I1(\mtime_compare[31]_i_3_n_0 ),
        .I2(\processor/wb_csr_address [6]),
        .I3(\processor/wb_csr_address [5]),
        .I4(\processor/wb_csr_address [0]),
        .I5(\mtvec[31]_i_2_n_0 ),
        .O(\mtvec[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \mtvec[31]_i_2 
       (.I0(\processor/wb_csr_address [3]),
        .I1(\processor/wb_csr_address [4]),
        .I2(\processor/wb_csr_address [1]),
        .I3(\processor/wb_csr_address [2]),
        .O(\mtvec[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[0]_i_1 
       (.I0(\processor/wb_csr_data [0]),
        .I1(mtvec[0]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(mtvec_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair100" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[10]_i_1 
       (.I0(\processor/wb_csr_data [10]),
        .I1(mtvec[10]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair123" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[11]_i_1 
       (.I0(\processor/wb_csr_data [11]),
        .I1(mtvec[11]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair124" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[12]_i_1 
       (.I0(\processor/wb_csr_data [12]),
        .I1(mtvec[12]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair125" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[13]_i_1 
       (.I0(\processor/wb_csr_data [13]),
        .I1(mtvec[13]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair96" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[14]_i_1 
       (.I0(\processor/wb_csr_data [14]),
        .I1(mtvec[14]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair126" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[15]_i_1 
       (.I0(\processor/wb_csr_data [15]),
        .I1(mtvec[15]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair126" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[16]_i_1 
       (.I0(\processor/wb_csr_data [16]),
        .I1(mtvec[16]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[16]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair128" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[17]_i_1 
       (.I0(\processor/wb_csr_data [17]),
        .I1(mtvec[17]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[17]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[18]_i_1 
       (.I0(\processor/wb_csr_data [18]),
        .I1(mtvec[18]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[18]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair129" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[19]_i_1 
       (.I0(\processor/wb_csr_data [19]),
        .I1(mtvec[19]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[19]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair92" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[1]_i_1 
       (.I0(\processor/wb_csr_data [1]),
        .I1(mtvec[1]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair130" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[20]_i_1 
       (.I0(\processor/wb_csr_data [20]),
        .I1(mtvec[20]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[20]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair131" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[21]_i_1 
       (.I0(\processor/wb_csr_data [21]),
        .I1(mtvec[21]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair132" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[22]_i_1 
       (.I0(\processor/wb_csr_data [22]),
        .I1(mtvec[22]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[22]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair132" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[23]_i_1 
       (.I0(\processor/wb_csr_data [23]),
        .I1(mtvec[23]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[23]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair131" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[24]_i_1 
       (.I0(\processor/wb_csr_data [24]),
        .I1(mtvec[24]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[24]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair130" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[25]_i_1 
       (.I0(\processor/wb_csr_data [25]),
        .I1(mtvec[25]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[25]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair129" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[26]_i_1 
       (.I0(\processor/wb_csr_data [26]),
        .I1(mtvec[26]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[26]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair128" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[27]_i_1 
       (.I0(\processor/wb_csr_data [27]),
        .I1(mtvec[27]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[27]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair125" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[28]_i_1 
       (.I0(\processor/wb_csr_data [28]),
        .I1(mtvec[28]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[28]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair124" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[29]_i_1 
       (.I0(\processor/wb_csr_data [29]),
        .I1(mtvec[29]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[29]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair92" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[2]_i_1 
       (.I0(\processor/wb_csr_data [2]),
        .I1(mtvec[2]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair123" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[30]_i_1 
       (.I0(\processor/wb_csr_data [30]),
        .I1(mtvec[30]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[30]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair122" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[31]_i_1 
       (.I0(\processor/wb_csr_data [31]),
        .I1(mtvec[31]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \mtvec_out[31]_i_2 
       (.I0(\mtvec_out[31]_i_3_n_0 ),
        .I1(\mtvec_out[31]_i_4_n_0 ),
        .I2(\processor/wb_csr_address [6]),
        .I3(\processor/wb_csr_address [7]),
        .I4(\processor/wb_csr_address [4]),
        .I5(\processor/wb_csr_address [5]),
        .O(\processor/csr_unit/mtvec_out1__6 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF1)) 
    \mtvec_out[31]_i_3 
       (.I0(\processor/wb_csr_write [0]),
        .I1(\processor/wb_csr_write [1]),
        .I2(\processor/wb_csr_address [2]),
        .I3(\processor/wb_csr_address [1]),
        .I4(\processor/wb_csr_address [11]),
        .I5(\processor/wb_csr_address [10]),
        .O(\mtvec_out[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2000)) 
    \mtvec_out[31]_i_4 
       (.I0(\processor/wb_csr_address [9]),
        .I1(\processor/wb_csr_address [3]),
        .I2(\processor/wb_csr_address [0]),
        .I3(\processor/wb_csr_address [8]),
        .O(\mtvec_out[31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair93" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[3]_i_1 
       (.I0(\processor/wb_csr_data [3]),
        .I1(mtvec[3]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair96" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[4]_i_1 
       (.I0(\processor/wb_csr_data [4]),
        .I1(mtvec[4]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair100" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[5]_i_1 
       (.I0(\processor/wb_csr_data [5]),
        .I1(mtvec[5]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair107" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[6]_i_1 
       (.I0(\processor/wb_csr_data [6]),
        .I1(mtvec[6]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair107" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[7]_i_1 
       (.I0(\processor/wb_csr_data [7]),
        .I1(mtvec[7]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair93" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[8]_i_1 
       (.I0(\processor/wb_csr_data [8]),
        .I1(mtvec[8]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair122" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \mtvec_out[9]_i_1 
       (.I0(\processor/wb_csr_data [9]),
        .I1(mtvec[9]),
        .I2(\processor/csr_unit/mtvec_out1__6 ),
        .O(\mtvec_out[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAA3F30)) 
    \pc[0]_i_1 
       (.I0(\processor/exception_target [0]),
        .I1(\pc[0]_i_3_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(pc[0]),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[0]_i_2 
       (.I0(\processor/mem_csr_data [0]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [0]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [0]),
        .O(\processor/exception_target [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCBFFFB)) 
    \pc[0]_i_3 
       (.I0(\csr_data_out[0]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[3]_i_4_n_7 ),
        .O(\pc[0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[10]_i_1 
       (.I0(\processor/exception_target [10]),
        .I1(\pc[10]_i_2_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[12]_i_4_n_6 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[10]_i_2 
       (.I0(\csr_data_out[10]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[11]_i_3_n_5 ),
        .O(\pc[10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[11]_i_1 
       (.I0(\processor/exception_target [11]),
        .I1(\pc[11]_i_2_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[12]_i_4_n_5 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[11]_i_2 
       (.I0(\csr_data_out[11]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[11]_i_3_n_4 ),
        .O(\pc[11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[11]_i_4 
       (.I0(\processor/execute/immediate [11]),
        .I1(\processor/execute/rs1_forwarded [11]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [11]),
        .O(\pc[11]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[11]_i_5 
       (.I0(\processor/execute/immediate [10]),
        .I1(\processor/execute/rs1_forwarded [10]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [10]),
        .O(\pc[11]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[11]_i_6 
       (.I0(\processor/execute/immediate [9]),
        .I1(\processor/execute/rs1_forwarded [9]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [9]),
        .O(\pc[11]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[11]_i_7 
       (.I0(\processor/execute/immediate [8]),
        .I1(\processor/execute/rs1_forwarded [8]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [8]),
        .O(\pc[11]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[12]_i_1 
       (.I0(\processor/exception_target [12]),
        .I1(\pc[12]_i_3_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[12]_i_4_n_4 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[12]_i_3 
       (.I0(\csr_data_out[12]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[15]_i_3_n_7 ),
        .O(\pc[12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[12]_i_5 
       (.I0(\processor/mem_csr_data [12]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [12]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [12]),
        .O(\processor/execute/mtvec_forwarded [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[12]_i_6 
       (.I0(\processor/mem_csr_data [11]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [11]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [11]),
        .O(\processor/execute/mtvec_forwarded [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[12]_i_7 
       (.I0(\processor/mem_csr_data [10]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [10]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [10]),
        .O(\processor/execute/mtvec_forwarded [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[12]_i_8 
       (.I0(\processor/mem_csr_data [9]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [9]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [9]),
        .O(\processor/execute/mtvec_forwarded [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[13]_i_1 
       (.I0(\processor/exception_target [13]),
        .I1(\pc[13]_i_2_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[16]_i_4_n_7 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[13]_i_2 
       (.I0(\csr_data_out[13]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[15]_i_3_n_6 ),
        .O(\pc[13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[14]_i_1 
       (.I0(\processor/exception_target [14]),
        .I1(\pc[14]_i_2_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[16]_i_4_n_6 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[14]_i_2 
       (.I0(\csr_data_out[14]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[15]_i_3_n_5 ),
        .O(\pc[14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[15]_i_1 
       (.I0(\processor/exception_target [15]),
        .I1(\pc[15]_i_2_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[16]_i_4_n_5 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[15]_i_2 
       (.I0(\csr_data_out[15]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[15]_i_3_n_4 ),
        .O(\pc[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[15]_i_4 
       (.I0(\processor/execute/immediate [15]),
        .I1(\processor/execute/rs1_forwarded [15]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [15]),
        .O(\pc[15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[15]_i_5 
       (.I0(\processor/execute/immediate [14]),
        .I1(\processor/execute/rs1_forwarded [14]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [14]),
        .O(\pc[15]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[15]_i_6 
       (.I0(\processor/execute/immediate [13]),
        .I1(\processor/execute/rs1_forwarded [13]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [13]),
        .O(\pc[15]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[15]_i_7 
       (.I0(\processor/execute/immediate [12]),
        .I1(\processor/execute/rs1_forwarded [12]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [12]),
        .O(\pc[15]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[16]_i_1 
       (.I0(\processor/exception_target [16]),
        .I1(\pc[16]_i_3_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[16]_i_4_n_4 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[16]_i_3 
       (.I0(\csr_data_out[16]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[19]_i_3_n_7 ),
        .O(\pc[16]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[16]_i_5 
       (.I0(\processor/mem_csr_data [16]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [16]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [16]),
        .O(\processor/execute/mtvec_forwarded [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[16]_i_6 
       (.I0(\processor/mem_csr_data [15]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [15]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [15]),
        .O(\processor/execute/mtvec_forwarded [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[16]_i_7 
       (.I0(\processor/mem_csr_data [14]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [14]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [14]),
        .O(\processor/execute/mtvec_forwarded [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[16]_i_8 
       (.I0(\processor/mem_csr_data [13]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [13]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [13]),
        .O(\processor/execute/mtvec_forwarded [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[17]_i_1 
       (.I0(\processor/exception_target [17]),
        .I1(\pc[17]_i_2_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[20]_i_4_n_7 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[17]_i_2 
       (.I0(\csr_data_out[17]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[19]_i_3_n_6 ),
        .O(\pc[17]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[18]_i_1 
       (.I0(\processor/exception_target [18]),
        .I1(\pc[18]_i_2_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[20]_i_4_n_6 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[18]_i_2 
       (.I0(\csr_data_out[18]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[19]_i_3_n_5 ),
        .O(\pc[18]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[19]_i_1 
       (.I0(\processor/exception_target [19]),
        .I1(\pc[19]_i_2_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[20]_i_4_n_5 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[19]_i_2 
       (.I0(\csr_data_out[19]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[19]_i_3_n_4 ),
        .O(\pc[19]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[19]_i_4 
       (.I0(\processor/execute/immediate [19]),
        .I1(\processor/execute/rs1_forwarded [19]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [19]),
        .O(\pc[19]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[19]_i_5 
       (.I0(\processor/execute/immediate [18]),
        .I1(\processor/execute/rs1_forwarded [18]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [18]),
        .O(\pc[19]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[19]_i_6 
       (.I0(\processor/execute/immediate [17]),
        .I1(\processor/execute/rs1_forwarded [17]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [17]),
        .O(\pc[19]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[19]_i_7 
       (.I0(\processor/execute/immediate [16]),
        .I1(\processor/execute/rs1_forwarded [16]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [16]),
        .O(\pc[19]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAA3F30)) 
    \pc[1]_i_1 
       (.I0(\processor/exception_target [1]),
        .I1(\pc[1]_i_3_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[4]_i_3_n_7 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[1]_i_2 
       (.I0(\processor/mem_csr_data [1]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [1]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [1]),
        .O(\processor/exception_target [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCBFFFB)) 
    \pc[1]_i_3 
       (.I0(\csr_data_out[1]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[3]_i_4_n_6 ),
        .O(\pc[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[20]_i_1 
       (.I0(\processor/exception_target [20]),
        .I1(\pc[20]_i_3_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[20]_i_4_n_4 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[20]_i_3 
       (.I0(\csr_data_out[20]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[23]_i_3_n_7 ),
        .O(\pc[20]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[20]_i_5 
       (.I0(\processor/mem_csr_data [20]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [20]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [20]),
        .O(\processor/execute/mtvec_forwarded [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[20]_i_6 
       (.I0(\processor/mem_csr_data [19]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [19]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [19]),
        .O(\processor/execute/mtvec_forwarded [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[20]_i_7 
       (.I0(\processor/mem_csr_data [18]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [18]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [18]),
        .O(\processor/execute/mtvec_forwarded [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[20]_i_8 
       (.I0(\processor/mem_csr_data [17]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [17]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [17]),
        .O(\processor/execute/mtvec_forwarded [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[21]_i_1 
       (.I0(\processor/exception_target [21]),
        .I1(\pc[21]_i_2_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[24]_i_4_n_7 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[21]_i_2 
       (.I0(\csr_data_out[21]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[23]_i_3_n_6 ),
        .O(\pc[21]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[22]_i_1 
       (.I0(\processor/exception_target [22]),
        .I1(\pc[22]_i_2_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[24]_i_4_n_6 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[22]_i_2 
       (.I0(\csr_data_out[22]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[23]_i_3_n_5 ),
        .O(\pc[22]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[23]_i_1 
       (.I0(\processor/exception_target [23]),
        .I1(\pc[23]_i_2_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[24]_i_4_n_5 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[23]_i_2 
       (.I0(\csr_data_out[23]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[23]_i_3_n_4 ),
        .O(\pc[23]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[23]_i_4 
       (.I0(\processor/execute/immediate [23]),
        .I1(\processor/execute/rs1_forwarded [23]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [23]),
        .O(\pc[23]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[23]_i_5 
       (.I0(\processor/execute/immediate [22]),
        .I1(\processor/execute/rs1_forwarded [22]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [22]),
        .O(\pc[23]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[23]_i_6 
       (.I0(\processor/execute/immediate [21]),
        .I1(\processor/execute/rs1_forwarded [21]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [21]),
        .O(\pc[23]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[23]_i_7 
       (.I0(\processor/execute/immediate [20]),
        .I1(\processor/execute/rs1_forwarded [20]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [20]),
        .O(\pc[23]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[24]_i_1 
       (.I0(\processor/exception_target [24]),
        .I1(\pc[24]_i_3_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[24]_i_4_n_4 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[24]_i_3 
       (.I0(\csr_data_out[24]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[27]_i_3_n_7 ),
        .O(\pc[24]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[24]_i_5 
       (.I0(\processor/mem_csr_data [24]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [24]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [24]),
        .O(\processor/execute/mtvec_forwarded [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[24]_i_6 
       (.I0(\processor/mem_csr_data [23]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [23]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [23]),
        .O(\processor/execute/mtvec_forwarded [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[24]_i_7 
       (.I0(\processor/mem_csr_data [22]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [22]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [22]),
        .O(\processor/execute/mtvec_forwarded [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[24]_i_8 
       (.I0(\processor/mem_csr_data [21]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [21]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [21]),
        .O(\processor/execute/mtvec_forwarded [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[25]_i_1 
       (.I0(\processor/exception_target [25]),
        .I1(\pc[25]_i_2_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[28]_i_4_n_7 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[25]_i_2 
       (.I0(\csr_data_out[25]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[27]_i_3_n_6 ),
        .O(\pc[25]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[26]_i_1 
       (.I0(\processor/exception_target [26]),
        .I1(\pc[26]_i_2_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[28]_i_4_n_6 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[26]_i_2 
       (.I0(\csr_data_out[26]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[27]_i_3_n_5 ),
        .O(\pc[26]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[27]_i_1 
       (.I0(\processor/exception_target [27]),
        .I1(\pc[27]_i_2_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[28]_i_4_n_5 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[27]_i_2 
       (.I0(\csr_data_out[27]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[27]_i_3_n_4 ),
        .O(\pc[27]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[27]_i_4 
       (.I0(\processor/execute/immediate [27]),
        .I1(\processor/execute/rs1_forwarded [27]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [27]),
        .O(\pc[27]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[27]_i_5 
       (.I0(\processor/execute/immediate [26]),
        .I1(\processor/execute/rs1_forwarded [26]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [26]),
        .O(\pc[27]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[27]_i_6 
       (.I0(\processor/execute/immediate [25]),
        .I1(\processor/execute/rs1_forwarded [25]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [25]),
        .O(\pc[27]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[27]_i_7 
       (.I0(\processor/execute/immediate [24]),
        .I1(\processor/execute/rs1_forwarded [24]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [24]),
        .O(\pc[27]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[28]_i_1 
       (.I0(\processor/exception_target [28]),
        .I1(\pc[28]_i_3_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[28]_i_4_n_4 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[28]_i_3 
       (.I0(\csr_data_out[28]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[31]_i_9_n_7 ),
        .O(\pc[28]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[28]_i_5 
       (.I0(\processor/mem_csr_data [28]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [28]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [28]),
        .O(\processor/execute/mtvec_forwarded [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[28]_i_6 
       (.I0(\processor/mem_csr_data [27]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [27]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [27]),
        .O(\processor/execute/mtvec_forwarded [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[28]_i_7 
       (.I0(\processor/mem_csr_data [26]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [26]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [26]),
        .O(\processor/execute/mtvec_forwarded [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[28]_i_8 
       (.I0(\processor/mem_csr_data [25]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [25]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [25]),
        .O(\processor/execute/mtvec_forwarded [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[29]_i_1 
       (.I0(\processor/exception_target [29]),
        .I1(\pc[29]_i_2_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[31]_i_5_n_7 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[29]_i_2 
       (.I0(\csr_data_out[29]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[31]_i_9_n_6 ),
        .O(\pc[29]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[2]_i_1 
       (.I0(\processor/exception_target [2]),
        .I1(\pc[2]_i_3_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[4]_i_3_n_6 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[2]_i_2 
       (.I0(\processor/mem_csr_data [2]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [2]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [2]),
        .O(\processor/exception_target [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[2]_i_3 
       (.I0(\csr_data_out[2]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[3]_i_4_n_5 ),
        .O(\pc[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[30]_i_1 
       (.I0(\processor/exception_target [30]),
        .I1(\pc[30]_i_2_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[31]_i_5_n_6 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[30]_i_2 
       (.I0(\csr_data_out[30]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[31]_i_9_n_5 ),
        .O(\pc[30]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00020000)) 
    \pc[31]_i_1 
       (.I0(imem_ack),
        .I1(\processor/fetch/cancel_fetch ),
        .I2(\mem_op[2]_i_5_n_0 ),
        .I3(\mem_op[2]_i_4_n_0 ),
        .I4(\processor/execute/exception_taken0 ),
        .O(\pc[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[31]_i_13 
       (.I0(\processor/execute/immediate [31]),
        .I1(\processor/execute/rs1_forwarded [31]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [31]),
        .O(\pc[31]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[31]_i_14 
       (.I0(\processor/execute/immediate [30]),
        .I1(\processor/execute/rs1_forwarded [30]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [30]),
        .O(\pc[31]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[31]_i_15 
       (.I0(\processor/execute/immediate [29]),
        .I1(\processor/execute/rs1_forwarded [29]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [29]),
        .O(\pc[31]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[31]_i_16 
       (.I0(\processor/execute/immediate [28]),
        .I1(\processor/execute/rs1_forwarded [28]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [28]),
        .O(\pc[31]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \pc[31]_i_1__0 
       (.I0(imem_ack),
        .I1(\processor/fetch/cancel_fetch ),
        .O(\pc[31]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[31]_i_2 
       (.I0(\processor/exception_target [31]),
        .I1(\pc[31]_i_4_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[31]_i_5_n_5 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[31]_i_4 
       (.I0(\csr_data_out[31]_i_4_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[31]_i_9_n_4 ),
        .O(\pc[31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[31]_i_6 
       (.I0(\processor/mem_csr_data [31]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [31]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [31]),
        .O(\processor/execute/mtvec_forwarded [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[31]_i_7 
       (.I0(\processor/mem_csr_data [30]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [30]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [30]),
        .O(\processor/execute/mtvec_forwarded [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[31]_i_8 
       (.I0(\processor/mem_csr_data [29]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [29]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [29]),
        .O(\processor/execute/mtvec_forwarded [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[3]_i_1 
       (.I0(\processor/exception_target [3]),
        .I1(\pc[3]_i_3_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[4]_i_3_n_5 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[3]_i_2 
       (.I0(\processor/mem_csr_data [3]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [3]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [3]),
        .O(\processor/exception_target [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[3]_i_3 
       (.I0(\csr_data_out[3]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[3]_i_4_n_4 ),
        .O(\pc[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[3]_i_5 
       (.I0(\processor/execute/immediate [3]),
        .I1(\processor/execute/rs1_forwarded [3]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [3]),
        .O(\pc[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[3]_i_6 
       (.I0(\processor/execute/immediate [2]),
        .I1(\processor/execute/rs1_forwarded [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [2]),
        .O(\pc[3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[3]_i_7 
       (.I0(\processor/execute/immediate [1]),
        .I1(\processor/execute/rs1_forwarded [1]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [1]),
        .O(\pc[3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[3]_i_8 
       (.I0(\processor/execute/immediate [0]),
        .I1(\processor/execute/rs1_forwarded [0]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [0]),
        .O(\pc[3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[4]_i_1 
       (.I0(\processor/exception_target [4]),
        .I1(\pc[4]_i_2_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[4]_i_3_n_4 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[4]_i_2 
       (.I0(\csr_data_out[4]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[7]_i_3_n_7 ),
        .O(\pc[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9AAA)) 
    \pc[4]_i_6 
       (.I0(pc[2]),
        .I1(\processor/fetch/cancel_fetch ),
        .I2(\processor/execute/exception_taken0 ),
        .I3(imem_ack),
        .O(\pc[4]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[5]_i_1 
       (.I0(\processor/exception_target [5]),
        .I1(\pc[5]_i_2_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[8]_i_3_n_7 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[5]_i_2 
       (.I0(\csr_data_out[5]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[7]_i_3_n_6 ),
        .O(\pc[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[6]_i_1 
       (.I0(\processor/exception_target [6]),
        .I1(\pc[6]_i_2_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[8]_i_3_n_6 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[6]_i_2 
       (.I0(\csr_data_out[6]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[7]_i_3_n_5 ),
        .O(\pc[6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[7]_i_1 
       (.I0(\processor/exception_target [7]),
        .I1(\pc[7]_i_2_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[8]_i_3_n_5 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[7]_i_2 
       (.I0(\csr_data_out[7]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[7]_i_3_n_4 ),
        .O(\pc[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[7]_i_4 
       (.I0(\processor/execute/immediate [7]),
        .I1(\processor/execute/rs1_forwarded [7]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [7]),
        .O(\pc[7]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[7]_i_5 
       (.I0(\processor/execute/immediate [6]),
        .I1(\processor/execute/rs1_forwarded [6]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [6]),
        .O(\pc[7]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[7]_i_6 
       (.I0(\processor/execute/immediate [5]),
        .I1(\processor/execute/rs1_forwarded [5]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [5]),
        .O(\pc[7]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h56A6)) 
    \pc[7]_i_7 
       (.I0(\processor/execute/immediate [4]),
        .I1(\processor/execute/rs1_forwarded [4]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_pc [4]),
        .O(\pc[7]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[8]_i_1 
       (.I0(\processor/exception_target [8]),
        .I1(\pc[8]_i_2_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[8]_i_3_n_4 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[8]_i_2 
       (.I0(\csr_data_out[8]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[11]_i_3_n_7 ),
        .O(\pc[8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    \pc[9]_i_1 
       (.I0(\processor/exception_target [9]),
        .I1(\pc[9]_i_2_n_0 ),
        .I2(\mem_op[2]_i_4_n_0 ),
        .I3(\pc_reg[12]_i_4_n_7 ),
        .I4(\mem_op[2]_i_5_n_0 ),
        .O(pc_next[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33340004)) 
    \pc[9]_i_2 
       (.I0(\csr_data_out[9]_i_3_n_0 ),
        .I1(\processor/ex_branch [2]),
        .I2(\processor/ex_branch [0]),
        .I3(\processor/ex_branch [1]),
        .I4(\pc_reg[11]_i_3_n_6 ),
        .O(\pc[9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \pc_reg[11]_i_3 
       (.CI(\pc_reg[7]_i_3_n_0 ),
        .CO(pc_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI(\processor/execute/immediate [11:8]),
        .O({\pc_reg[11]_i_3_n_4 ,\pc_reg[11]_i_3_n_5 ,\pc_reg[11]_i_3_n_6 ,\pc_reg[11]_i_3_n_7 }),
        .S({\pc[11]_i_4_n_0 ,\pc[11]_i_5_n_0 ,\pc[11]_i_6_n_0 ,\pc[11]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \pc_reg[12]_i_2 
       (.CI(tag_memory_reg_0_63_0_2_i_8_n_0),
        .CO({\pc_reg[12]_i_2_n_0 ,\pc_reg[12]_i_2_n_1 ,\pc_reg[12]_i_2_n_2 ,\pc_reg[12]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\processor/exception_target [12:9]),
        .S(\processor/execute/mtvec_forwarded [12:9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \pc_reg[12]_i_4 
       (.CI(\pc_reg[8]_i_3_n_0 ),
        .CO({\pc_reg[12]_i_4_n_0 ,\pc_reg[12]_i_4_n_1 ,\pc_reg[12]_i_4_n_2 ,\pc_reg[12]_i_4_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\pc_reg[12]_i_4_n_4 ,\pc_reg[12]_i_4_n_5 ,\pc_reg[12]_i_4_n_6 ,\pc_reg[12]_i_4_n_7 }),
        .S(pc[12:9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \pc_reg[15]_i_3 
       (.CI(pc_reg[3]),
        .CO({\pc_reg[15]_i_3_n_0 ,\pc_reg[15]_i_3_n_1 ,\pc_reg[15]_i_3_n_2 ,\pc_reg[15]_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\processor/execute/immediate [15:12]),
        .O({\pc_reg[15]_i_3_n_4 ,\pc_reg[15]_i_3_n_5 ,\pc_reg[15]_i_3_n_6 ,\pc_reg[15]_i_3_n_7 }),
        .S({\pc[15]_i_4_n_0 ,\pc[15]_i_5_n_0 ,\pc[15]_i_6_n_0 ,\pc[15]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \pc_reg[16]_i_2 
       (.CI(\pc_reg[12]_i_2_n_0 ),
        .CO({\pc_reg[16]_i_2_n_0 ,\pc_reg[16]_i_2_n_1 ,\pc_reg[16]_i_2_n_2 ,\pc_reg[16]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\processor/exception_target [16:13]),
        .S(\processor/execute/mtvec_forwarded [16:13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \pc_reg[16]_i_4 
       (.CI(\pc_reg[12]_i_4_n_0 ),
        .CO({\pc_reg[16]_i_4_n_0 ,\pc_reg[16]_i_4_n_1 ,\pc_reg[16]_i_4_n_2 ,\pc_reg[16]_i_4_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\pc_reg[16]_i_4_n_4 ,\pc_reg[16]_i_4_n_5 ,\pc_reg[16]_i_4_n_6 ,\pc_reg[16]_i_4_n_7 }),
        .S(pc[16:13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \pc_reg[19]_i_3 
       (.CI(\pc_reg[15]_i_3_n_0 ),
        .CO({\pc_reg[19]_i_3_n_0 ,\pc_reg[19]_i_3_n_1 ,\pc_reg[19]_i_3_n_2 ,\pc_reg[19]_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\processor/execute/immediate [19:16]),
        .O({\pc_reg[19]_i_3_n_4 ,\pc_reg[19]_i_3_n_5 ,\pc_reg[19]_i_3_n_6 ,\pc_reg[19]_i_3_n_7 }),
        .S({\pc[19]_i_4_n_0 ,\pc[19]_i_5_n_0 ,\pc[19]_i_6_n_0 ,\pc[19]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \pc_reg[20]_i_2 
       (.CI(\pc_reg[16]_i_2_n_0 ),
        .CO({\pc_reg[20]_i_2_n_0 ,\pc_reg[20]_i_2_n_1 ,\pc_reg[20]_i_2_n_2 ,\pc_reg[20]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\processor/exception_target [20:17]),
        .S(\processor/execute/mtvec_forwarded [20:17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \pc_reg[20]_i_4 
       (.CI(\pc_reg[16]_i_4_n_0 ),
        .CO({\pc_reg[20]_i_4_n_0 ,\pc_reg[20]_i_4_n_1 ,\pc_reg[20]_i_4_n_2 ,\pc_reg[20]_i_4_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\pc_reg[20]_i_4_n_4 ,\pc_reg[20]_i_4_n_5 ,\pc_reg[20]_i_4_n_6 ,\pc_reg[20]_i_4_n_7 }),
        .S(pc[20:17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \pc_reg[23]_i_3 
       (.CI(\pc_reg[19]_i_3_n_0 ),
        .CO({\pc_reg[23]_i_3_n_0 ,\pc_reg[23]_i_3_n_1 ,\pc_reg[23]_i_3_n_2 ,\pc_reg[23]_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\processor/execute/immediate [23:20]),
        .O({\pc_reg[23]_i_3_n_4 ,\pc_reg[23]_i_3_n_5 ,\pc_reg[23]_i_3_n_6 ,\pc_reg[23]_i_3_n_7 }),
        .S({\pc[23]_i_4_n_0 ,\pc[23]_i_5_n_0 ,\pc[23]_i_6_n_0 ,\pc[23]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \pc_reg[24]_i_2 
       (.CI(\pc_reg[20]_i_2_n_0 ),
        .CO({\pc_reg[24]_i_2_n_0 ,\pc_reg[24]_i_2_n_1 ,\pc_reg[24]_i_2_n_2 ,\pc_reg[24]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\processor/exception_target [24:21]),
        .S(\processor/execute/mtvec_forwarded [24:21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \pc_reg[24]_i_4 
       (.CI(\pc_reg[20]_i_4_n_0 ),
        .CO({\pc_reg[24]_i_4_n_0 ,\pc_reg[24]_i_4_n_1 ,\pc_reg[24]_i_4_n_2 ,\pc_reg[24]_i_4_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\pc_reg[24]_i_4_n_4 ,\pc_reg[24]_i_4_n_5 ,\pc_reg[24]_i_4_n_6 ,\pc_reg[24]_i_4_n_7 }),
        .S(pc[24:21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \pc_reg[27]_i_3 
       (.CI(\pc_reg[23]_i_3_n_0 ),
        .CO({\pc_reg[27]_i_3_n_0 ,\pc_reg[27]_i_3_n_1 ,\pc_reg[27]_i_3_n_2 ,\pc_reg[27]_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\processor/execute/immediate [27:24]),
        .O({\pc_reg[27]_i_3_n_4 ,\pc_reg[27]_i_3_n_5 ,\pc_reg[27]_i_3_n_6 ,\pc_reg[27]_i_3_n_7 }),
        .S({\pc[27]_i_4_n_0 ,\pc[27]_i_5_n_0 ,\pc[27]_i_6_n_0 ,\pc[27]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \pc_reg[28]_i_2 
       (.CI(\pc_reg[24]_i_2_n_0 ),
        .CO({\pc_reg[28]_i_2_n_0 ,\pc_reg[28]_i_2_n_1 ,\pc_reg[28]_i_2_n_2 ,\pc_reg[28]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\processor/exception_target [28:25]),
        .S(\processor/execute/mtvec_forwarded [28:25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \pc_reg[28]_i_4 
       (.CI(\pc_reg[24]_i_4_n_0 ),
        .CO({\pc_reg[28]_i_4_n_0 ,\pc_reg[28]_i_4_n_1 ,\pc_reg[28]_i_4_n_2 ,\pc_reg[28]_i_4_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\pc_reg[28]_i_4_n_4 ,\pc_reg[28]_i_4_n_5 ,\pc_reg[28]_i_4_n_6 ,\pc_reg[28]_i_4_n_7 }),
        .S(pc[28:25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \pc_reg[31]_i_3 
       (.CI(\pc_reg[28]_i_2_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\pc_reg[31]_i_3_n_4 ,\processor/exception_target [31:29]}),
        .S({\<const0>__0__0 ,\processor/execute/mtvec_forwarded [31:29]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \pc_reg[31]_i_5 
       (.CI(\pc_reg[28]_i_4_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\pc_reg[31]_i_5_n_4 ,\pc_reg[31]_i_5_n_5 ,\pc_reg[31]_i_5_n_6 ,\pc_reg[31]_i_5_n_7 }),
        .S({\<const0>__0__0 ,pc[31:29]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \pc_reg[31]_i_9 
       (.CI(\pc_reg[27]_i_3_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\processor/execute/immediate [30:28]}),
        .O({\pc_reg[31]_i_9_n_4 ,\pc_reg[31]_i_9_n_5 ,\pc_reg[31]_i_9_n_6 ,\pc_reg[31]_i_9_n_7 }),
        .S({\pc[31]_i_13_n_0 ,\pc[31]_i_14_n_0 ,\pc[31]_i_15_n_0 ,\pc[31]_i_16_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \pc_reg[3]_i_4 
       (.CI(\<const0>__0__0 ),
        .CO({\pc_reg[3]_i_4_n_0 ,\pc_reg[3]_i_4_n_1 ,\pc_reg[3]_i_4_n_2 ,\pc_reg[3]_i_4_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\processor/execute/immediate [3:0]),
        .O({\pc_reg[3]_i_4_n_4 ,\pc_reg[3]_i_4_n_5 ,\pc_reg[3]_i_4_n_6 ,\pc_reg[3]_i_4_n_7 }),
        .S({\pc[3]_i_5_n_0 ,\pc[3]_i_6_n_0 ,\pc[3]_i_7_n_0 ,\pc[3]_i_8_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \pc_reg[4]_i_3 
       (.CI(\<const0>__0__0 ),
        .CO({\pc_reg[4]_i_3_n_0 ,\pc_reg[4]_i_3_n_1 ,\pc_reg[4]_i_3_n_2 ,\pc_reg[4]_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,pc[2],\<const0>__0__0 }),
        .O({\pc_reg[4]_i_3_n_4 ,\pc_reg[4]_i_3_n_5 ,\pc_reg[4]_i_3_n_6 ,\pc_reg[4]_i_3_n_7 }),
        .S({pc[4:3],\pc[4]_i_6_n_0 ,pc[1]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \pc_reg[7]_i_3 
       (.CI(\pc_reg[3]_i_4_n_0 ),
        .CO({\pc_reg[7]_i_3_n_0 ,\pc_reg[7]_i_3_n_1 ,\pc_reg[7]_i_3_n_2 ,\pc_reg[7]_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\processor/execute/immediate [7:4]),
        .O({\pc_reg[7]_i_3_n_4 ,\pc_reg[7]_i_3_n_5 ,\pc_reg[7]_i_3_n_6 ,\pc_reg[7]_i_3_n_7 }),
        .S({\pc[7]_i_4_n_0 ,\pc[7]_i_5_n_0 ,\pc[7]_i_6_n_0 ,\pc[7]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \pc_reg[8]_i_3 
       (.CI(\pc_reg[4]_i_3_n_0 ),
        .CO({\pc_reg[8]_i_3_n_0 ,\pc_reg[8]_i_3_n_1 ,\pc_reg[8]_i_3_n_2 ,\pc_reg[8]_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\pc_reg[8]_i_3_n_4 ,\pc_reg[8]_i_3_n_5 ,\pc_reg[8]_i_3_n_6 ,\pc_reg[8]_i_3_n_7 }),
        .S(pc[8:5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_read_address_p_reg[0] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/decode/csr_addr__40 [0]),
        .Q(csr_read_address_p[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_read_address_p_reg[10] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_immediate [10]),
        .Q(csr_read_address_p[10]),
        .R(\csr_read_address_p[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_read_address_p_reg[11] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_immediate [11]),
        .Q(csr_read_address_p[11]),
        .R(\csr_read_address_p[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_read_address_p_reg[1] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_immediate [1]),
        .Q(csr_read_address_p[1]),
        .R(\csr_read_address_p[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_read_address_p_reg[2] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_immediate [2]),
        .Q(csr_read_address_p[2]),
        .R(\csr_read_address_p[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_read_address_p_reg[3] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_immediate [3]),
        .Q(csr_read_address_p[3]),
        .R(\csr_read_address_p[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_read_address_p_reg[4] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_immediate [4]),
        .Q(csr_read_address_p[4]),
        .R(\csr_read_address_p[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_read_address_p_reg[5] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_immediate [5]),
        .Q(csr_read_address_p[5]),
        .R(\csr_read_address_p[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_read_address_p_reg[6] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/decode/csr_addr__40 [6]),
        .Q(csr_read_address_p[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_read_address_p_reg[7] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_immediate [7]),
        .Q(csr_read_address_p[7]),
        .R(\csr_read_address_p[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_read_address_p_reg[8] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/decode/csr_addr__40 [8]),
        .Q(csr_read_address_p[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_read_address_p_reg[9] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/decode/csr_addr__40 [9]),
        .Q(csr_read_address_p[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[0] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[0]_i_1_n_7 ),
        .Q(\processor/csr_unit/counter_mtime_reg [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[10] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[8]_i_1_n_5 ),
        .Q(\processor/csr_unit/counter_mtime_reg [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[11] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[8]_i_1_n_4 ),
        .Q(\processor/csr_unit/counter_mtime_reg [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[12] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[12]_i_1_n_7 ),
        .Q(\processor/csr_unit/counter_mtime_reg [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[13] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[12]_i_1_n_6 ),
        .Q(\processor/csr_unit/counter_mtime_reg [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[14] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[12]_i_1_n_5 ),
        .Q(\processor/csr_unit/counter_mtime_reg [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[15] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[12]_i_1_n_4 ),
        .Q(\processor/csr_unit/counter_mtime_reg [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[16] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[16]_i_1_n_7 ),
        .Q(\processor/csr_unit/counter_mtime_reg [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[17] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[16]_i_1_n_6 ),
        .Q(\processor/csr_unit/counter_mtime_reg [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[18] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[16]_i_1_n_5 ),
        .Q(\processor/csr_unit/counter_mtime_reg [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[19] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[16]_i_1_n_4 ),
        .Q(\processor/csr_unit/counter_mtime_reg [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[1] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[0]_i_1_n_6 ),
        .Q(\processor/csr_unit/counter_mtime_reg [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[20] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[20]_i_1_n_7 ),
        .Q(\processor/csr_unit/counter_mtime_reg [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[21] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[20]_i_1_n_6 ),
        .Q(\processor/csr_unit/counter_mtime_reg [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[22] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[20]_i_1_n_5 ),
        .Q(\processor/csr_unit/counter_mtime_reg [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[23] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[20]_i_1_n_4 ),
        .Q(\processor/csr_unit/counter_mtime_reg [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[24] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[24]_i_1_n_7 ),
        .Q(\processor/csr_unit/counter_mtime_reg [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[25] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[24]_i_1_n_6 ),
        .Q(\processor/csr_unit/counter_mtime_reg [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[26] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[24]_i_1_n_5 ),
        .Q(\processor/csr_unit/counter_mtime_reg [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[27] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[24]_i_1_n_4 ),
        .Q(\processor/csr_unit/counter_mtime_reg [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[28] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[28]_i_1_n_7 ),
        .Q(\processor/csr_unit/counter_mtime_reg [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[29] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[28]_i_1_n_6 ),
        .Q(\processor/csr_unit/counter_mtime_reg [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[2] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[0]_i_1_n_5 ),
        .Q(\processor/csr_unit/counter_mtime_reg [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[30] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[28]_i_1_n_5 ),
        .Q(\processor/csr_unit/counter_mtime_reg [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[31] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[28]_i_1_n_4 ),
        .Q(\processor/csr_unit/counter_mtime_reg [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[3] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[0]_i_1_n_4 ),
        .Q(\processor/csr_unit/counter_mtime_reg [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[4] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[4]_i_1_n_7 ),
        .Q(\processor/csr_unit/counter_mtime_reg [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[5] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[4]_i_1_n_6 ),
        .Q(\processor/csr_unit/counter_mtime_reg [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[6] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[4]_i_1_n_5 ),
        .Q(\processor/csr_unit/counter_mtime_reg [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[7] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[4]_i_1_n_4 ),
        .Q(\processor/csr_unit/counter_mtime_reg [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[8] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[8]_i_1_n_7 ),
        .Q(\processor/csr_unit/counter_mtime_reg [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \processor/csr_unit/counter_mtime_reg[9] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(\counter_mtime_reg[8]_i_1_n_6 ),
        .Q(\processor/csr_unit/counter_mtime_reg [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[0]_i_1__0_n_7 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_ ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[8]_i_1__0_n_5 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[10] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[8]_i_1__0_n_4 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[11] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[12]_i_1__0_n_7 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[12] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[12]_i_1__0_n_6 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[13] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[12]_i_1__0_n_5 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[14] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[12]_i_1__0_n_4 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[15] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[16]_i_1__0_n_7 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[16] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[16]_i_1__0_n_6 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[17] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[16]_i_1__0_n_5 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[18] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[16]_i_1__0_n_4 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[19] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[0]_i_1__0_n_6 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[1] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[20]_i_1__0_n_7 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[20] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[20]_i_1__0_n_6 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[21] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[20]_i_1__0_n_5 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[22] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[20]_i_1__0_n_4 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[23] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[24]_i_1__0_n_7 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[24] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[24]_i_1__0_n_6 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[25] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[24]_i_1__0_n_5 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[26] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[24]_i_1__0_n_4 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[27] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[28]_i_1__0_n_7 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[28] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[28]_i_1__0_n_6 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[29] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[0]_i_1__0_n_5 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[2] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[28]_i_1__0_n_5 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[30] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[28]_i_1__0_n_4 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[31] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[32]_i_1__0_n_7 ),
        .Q(data14[0]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[32]_i_1__0_n_6 ),
        .Q(data14[1]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[32]_i_1__0_n_5 ),
        .Q(data14[2]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[32]_i_1__0_n_4 ),
        .Q(data14[3]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[36]_i_1__0_n_7 ),
        .Q(data14[4]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[36]_i_1__0_n_6 ),
        .Q(data14[5]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[36]_i_1__0_n_5 ),
        .Q(data14[6]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[36]_i_1__0_n_4 ),
        .Q(data14[7]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[0]_i_1__0_n_4 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[3] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[40]_i_1__0_n_7 ),
        .Q(data14[8]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[40]_i_1__0_n_6 ),
        .Q(data14[9]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[40]_i_1__0_n_5 ),
        .Q(data14[10]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[40]_i_1__0_n_4 ),
        .Q(data14[11]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[44]_i_1__0_n_7 ),
        .Q(data14[12]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[44]_i_1__0_n_6 ),
        .Q(data14[13]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[44]_i_1__0_n_5 ),
        .Q(data14[14]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[44]_i_1__0_n_4 ),
        .Q(data14[15]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[48]_i_1__0_n_7 ),
        .Q(data14[16]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[48]_i_1__0_n_6 ),
        .Q(data14[17]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[4]_i_1__0_n_7 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[4] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[48]_i_1__0_n_5 ),
        .Q(data14[18]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[48]_i_1__0_n_4 ),
        .Q(data14[19]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[52]_i_1__0_n_7 ),
        .Q(data14[20]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[52]_i_1__0_n_6 ),
        .Q(data14[21]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[52]_i_1__0_n_5 ),
        .Q(data14[22]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[52]_i_1__0_n_4 ),
        .Q(data14[23]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[56]_i_1__0_n_7 ),
        .Q(data14[24]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[56]_i_1__0_n_6 ),
        .Q(data14[25]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[56]_i_1__0_n_5 ),
        .Q(data14[26]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[56]_i_1__0_n_4 ),
        .Q(data14[27]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[4]_i_1__0_n_6 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[5] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[60]_i_1__0_n_7 ),
        .Q(data14[28]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[60]_i_1__0_n_6 ),
        .Q(data14[29]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[60]_i_1__0_n_5 ),
        .Q(data14[30]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[60]_i_1__0_n_4 ),
        .Q(data14[31]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[4]_i_1__0_n_5 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[6] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[4]_i_1__0_n_4 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[7] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[8]_i_1__0_n_7 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[8] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/cycle_counter/current_count_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[8]_i_1__0_n_6 ),
        .Q(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[9] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[0] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[0]),
        .Q(fromhost[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[10] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[10]),
        .Q(fromhost[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[11] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[11]),
        .Q(fromhost[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[12] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[12]),
        .Q(fromhost[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[13] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[13]),
        .Q(fromhost[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[14] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[14]),
        .Q(fromhost[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[15] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[15]),
        .Q(fromhost[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[16] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[16]),
        .Q(fromhost[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[17] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[17]),
        .Q(fromhost[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[18] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[18]),
        .Q(fromhost[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[19] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[19]),
        .Q(fromhost[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[1] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[1]),
        .Q(fromhost[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[20] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[20]),
        .Q(fromhost[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[21] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[21]),
        .Q(fromhost[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[22] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[22]),
        .Q(fromhost[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[23] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[23]),
        .Q(fromhost[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[24] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[24]),
        .Q(fromhost[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[25] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[25]),
        .Q(fromhost[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[26] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[26]),
        .Q(fromhost[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[27] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[27]),
        .Q(fromhost[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[28] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[28]),
        .Q(fromhost[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[29] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[29]),
        .Q(fromhost[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[2] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[2]),
        .Q(fromhost[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[30] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[30]),
        .Q(fromhost[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[31] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[31]),
        .Q(fromhost[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[3] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[3]),
        .Q(fromhost[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[4] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[4]),
        .Q(fromhost[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[5] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[5]),
        .Q(fromhost[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[6] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[6]),
        .Q(fromhost[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[7] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[7]),
        .Q(fromhost[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[8] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[8]),
        .Q(fromhost[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/fromhost_reg[9] 
       (.C(clk),
        .CE(fromhost_updated),
        .D(fromhost_data[9]),
        .Q(fromhost[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/ie1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(ie1_i_1_n_0),
        .Q(\processor/ie1 ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/ie_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(ie_i_1_n_0),
        .Q(\processor/ie ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[0] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[0]_i_1__1_n_7 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_ ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[10] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[8]_i_1__1_n_5 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[10] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[11] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[8]_i_1__1_n_4 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[11] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[12] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[12]_i_1__1_n_7 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[12] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[13] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[12]_i_1__1_n_6 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[13] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[14] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[12]_i_1__1_n_5 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[14] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[15] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[12]_i_1__1_n_4 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[15] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[16] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[16]_i_1__1_n_7 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[16] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[17] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[16]_i_1__1_n_6 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[17] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[18] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[16]_i_1__1_n_5 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[18] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[19] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[16]_i_1__1_n_4 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[19] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[1] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[0]_i_1__1_n_6 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[1] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[20] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[20]_i_1__1_n_7 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[20] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[21] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[20]_i_1__1_n_6 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[21] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[22] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[20]_i_1__1_n_5 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[22] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[23] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[20]_i_1__1_n_4 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[23] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[24] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[24]_i_1__1_n_7 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[24] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[25] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[24]_i_1__1_n_6 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[25] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[26] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[24]_i_1__1_n_5 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[26] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[27] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[24]_i_1__1_n_4 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[27] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[28] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[28]_i_1__1_n_7 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[28] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[29] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[28]_i_1__1_n_6 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[29] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[2] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[0]_i_1__1_n_5 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[2] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[30] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[28]_i_1__1_n_5 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[30] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[31] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[28]_i_1__1_n_4 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[31] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[32] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[32]_i_1__1_n_7 ),
        .Q(data16[0]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[33] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[32]_i_1__1_n_6 ),
        .Q(data16[1]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[34] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[32]_i_1__1_n_5 ),
        .Q(data16[2]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[35] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[32]_i_1__1_n_4 ),
        .Q(data16[3]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[36] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[36]_i_1__1_n_7 ),
        .Q(data16[4]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[37] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[36]_i_1__1_n_6 ),
        .Q(data16[5]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[38] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[36]_i_1__1_n_5 ),
        .Q(data16[6]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[39] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[36]_i_1__1_n_4 ),
        .Q(data16[7]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[3] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[0]_i_1__1_n_4 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[3] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[40] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[40]_i_1__1_n_7 ),
        .Q(data16[8]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[41] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[40]_i_1__1_n_6 ),
        .Q(data16[9]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[42] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[40]_i_1__1_n_5 ),
        .Q(data16[10]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[43] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[40]_i_1__1_n_4 ),
        .Q(data16[11]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[44] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[44]_i_1__1_n_7 ),
        .Q(data16[12]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[45] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[44]_i_1__1_n_6 ),
        .Q(data16[13]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[46] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[44]_i_1__1_n_5 ),
        .Q(data16[14]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[47] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[44]_i_1__1_n_4 ),
        .Q(data16[15]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[48] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[48]_i_1__1_n_7 ),
        .Q(data16[16]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[49] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[48]_i_1__1_n_6 ),
        .Q(data16[17]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[4] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[4]_i_1__1_n_7 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[4] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[50] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[48]_i_1__1_n_5 ),
        .Q(data16[18]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[51] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[48]_i_1__1_n_4 ),
        .Q(data16[19]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[52] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[52]_i_1__1_n_7 ),
        .Q(data16[20]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[53] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[52]_i_1__1_n_6 ),
        .Q(data16[21]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[54] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[52]_i_1__1_n_5 ),
        .Q(data16[22]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[55] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[52]_i_1__1_n_4 ),
        .Q(data16[23]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[56] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[56]_i_1__1_n_7 ),
        .Q(data16[24]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[57] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[56]_i_1__1_n_6 ),
        .Q(data16[25]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[58] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[56]_i_1__1_n_5 ),
        .Q(data16[26]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[59] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[56]_i_1__1_n_4 ),
        .Q(data16[27]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[5] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[4]_i_1__1_n_6 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[5] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[60] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[60]_i_1__1_n_7 ),
        .Q(data16[28]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[61] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[60]_i_1__1_n_6 ),
        .Q(data16[29]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[62] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[60]_i_1__1_n_5 ),
        .Q(data16[30]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[63] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[60]_i_1__1_n_4 ),
        .Q(data16[31]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[6] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[4]_i_1__1_n_5 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[6] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[7] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[4]_i_1__1_n_4 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[7] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[8] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[8]_i_1__1_n_7 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[8] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/instret_counter/current_count_reg[9] 
       (.C(clk),
        .CE(\processor/writeback/count_instr_out_reg_n_0 ),
        .D(\current_count_reg[8]_i_1__1_n_6 ),
        .Q(\processor/csr_unit/instret_counter/current_count_reg_n_0_[9] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[0] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [0]),
        .Q(mbadaddr[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[10] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [10]),
        .Q(mbadaddr[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[11] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [11]),
        .Q(mbadaddr[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[12] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [12]),
        .Q(mbadaddr[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[13] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [13]),
        .Q(mbadaddr[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[14] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [14]),
        .Q(mbadaddr[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[15] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [15]),
        .Q(mbadaddr[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[16] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [16]),
        .Q(mbadaddr[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[17] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [17]),
        .Q(mbadaddr[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[18] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [18]),
        .Q(mbadaddr[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[19] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [19]),
        .Q(mbadaddr[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[1] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [1]),
        .Q(mbadaddr[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[20] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [20]),
        .Q(mbadaddr[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[21] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [21]),
        .Q(mbadaddr[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[22] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [22]),
        .Q(mbadaddr[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[23] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [23]),
        .Q(mbadaddr[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[24] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [24]),
        .Q(mbadaddr[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[25] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [25]),
        .Q(mbadaddr[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[26] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [26]),
        .Q(mbadaddr[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[27] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [27]),
        .Q(mbadaddr[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[28] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [28]),
        .Q(mbadaddr[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[29] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [29]),
        .Q(mbadaddr[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[2] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [2]),
        .Q(mbadaddr[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[30] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [30]),
        .Q(mbadaddr[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[31] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [31]),
        .Q(mbadaddr[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[3] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [3]),
        .Q(mbadaddr[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[4] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [4]),
        .Q(mbadaddr[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[5] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [5]),
        .Q(mbadaddr[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[6] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [6]),
        .Q(mbadaddr[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[7] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [7]),
        .Q(mbadaddr[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[8] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [8]),
        .Q(mbadaddr[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mbadaddr_reg[9] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[badaddr] [9]),
        .Q(mbadaddr[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mcause_reg[0] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[cause] [0]),
        .Q(data8[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mcause_reg[1] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[cause] [1]),
        .Q(data8[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mcause_reg[2] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[cause] [2]),
        .Q(data8[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mcause_reg[3] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[cause] [3]),
        .Q(data8[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mcause_reg[4] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[cause] [4]),
        .Q(data8[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mcause_reg[5] 
       (.C(clk),
        .CE(\mbadaddr[31]_i_1_n_0 ),
        .D(\processor/wb_exception_context[cause] [5]),
        .Q(data8[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[0] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [0]),
        .Q(mepc[0]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[10] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [10]),
        .Q(mepc[10]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[11] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [11]),
        .Q(mepc[11]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[12] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [12]),
        .Q(mepc[12]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[13] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [13]),
        .Q(mepc[13]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[14] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [14]),
        .Q(mepc[14]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[15] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [15]),
        .Q(mepc[15]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[16] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [16]),
        .Q(mepc[16]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[17] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [17]),
        .Q(mepc[17]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[18] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [18]),
        .Q(mepc[18]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[19] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [19]),
        .Q(mepc[19]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[1] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [1]),
        .Q(mepc[1]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[20] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [20]),
        .Q(mepc[20]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[21] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [21]),
        .Q(mepc[21]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[22] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [22]),
        .Q(mepc[22]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[23] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [23]),
        .Q(mepc[23]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[24] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [24]),
        .Q(mepc[24]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[25] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [25]),
        .Q(mepc[25]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[26] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [26]),
        .Q(mepc[26]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[27] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [27]),
        .Q(mepc[27]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[28] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [28]),
        .Q(mepc[28]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[29] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [29]),
        .Q(mepc[29]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[2] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [2]),
        .Q(mepc[2]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[30] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [30]),
        .Q(mepc[30]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[31] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [31]),
        .Q(mepc[31]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[3] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [3]),
        .Q(mepc[3]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[4] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [4]),
        .Q(mepc[4]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[5] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [5]),
        .Q(mepc[5]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[6] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [6]),
        .Q(mepc[6]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[7] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [7]),
        .Q(mepc[7]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[8] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [8]),
        .Q(mepc[8]),
        .S(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mepc_reg[9] 
       (.C(clk),
        .CE(\mepc[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [9]),
        .Q(mepc[9]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[0] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [0]),
        .Q(\processor/mie [0]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[10] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [10]),
        .Q(\processor/mie [10]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[11] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [11]),
        .Q(\processor/mie [11]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[12] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [12]),
        .Q(\processor/mie [12]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[13] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [13]),
        .Q(\processor/mie [13]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[14] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [14]),
        .Q(\processor/mie [14]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[15] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [15]),
        .Q(\processor/mie [15]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[16] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [16]),
        .Q(\processor/mie [16]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[17] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [17]),
        .Q(\processor/mie [17]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[18] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [18]),
        .Q(\processor/mie [18]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[19] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [19]),
        .Q(\processor/mie [19]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[1] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [1]),
        .Q(\processor/mie [1]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[20] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [20]),
        .Q(\processor/mie [20]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[21] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [21]),
        .Q(\processor/mie [21]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[22] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [22]),
        .Q(\processor/mie [22]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[23] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [23]),
        .Q(\processor/mie [23]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[24] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [24]),
        .Q(\processor/mie [24]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[25] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [25]),
        .Q(\processor/mie [25]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[26] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [26]),
        .Q(\processor/mie [26]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[27] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [27]),
        .Q(\processor/mie [27]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[28] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [28]),
        .Q(\processor/mie [28]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[29] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [29]),
        .Q(\processor/mie [29]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[2] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [2]),
        .Q(\processor/mie [2]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[30] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [30]),
        .Q(\processor/mie [30]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[31] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [31]),
        .Q(\processor/mie [31]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[3] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [3]),
        .Q(\processor/mie [3]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[4] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [4]),
        .Q(\processor/mie [4]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[5] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [5]),
        .Q(\processor/mie [5]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[6] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [6]),
        .Q(\processor/mie [6]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[7] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [7]),
        .Q(\processor/mie [7]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[8] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [8]),
        .Q(\processor/mie [8]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mie_reg[9] 
       (.C(clk),
        .CE(mie),
        .D(\processor/wb_csr_data [9]),
        .Q(\processor/mie [9]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[0] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [0]),
        .Q(mscratch[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[10] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [10]),
        .Q(mscratch[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[11] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [11]),
        .Q(mscratch[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[12] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [12]),
        .Q(mscratch[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[13] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [13]),
        .Q(mscratch[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[14] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [14]),
        .Q(mscratch[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[15] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [15]),
        .Q(mscratch[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[16] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [16]),
        .Q(mscratch[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[17] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [17]),
        .Q(mscratch[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[18] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [18]),
        .Q(mscratch[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[19] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [19]),
        .Q(mscratch[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[1] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [1]),
        .Q(mscratch[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[20] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [20]),
        .Q(mscratch[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[21] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [21]),
        .Q(mscratch[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[22] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [22]),
        .Q(mscratch[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[23] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [23]),
        .Q(mscratch[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[24] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [24]),
        .Q(mscratch[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[25] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [25]),
        .Q(mscratch[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[26] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [26]),
        .Q(mscratch[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[27] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [27]),
        .Q(mscratch[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[28] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [28]),
        .Q(mscratch[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[29] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [29]),
        .Q(mscratch[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[2] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [2]),
        .Q(mscratch[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[30] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [30]),
        .Q(mscratch[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[31] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [31]),
        .Q(mscratch[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[3] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [3]),
        .Q(mscratch[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[4] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [4]),
        .Q(mscratch[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[5] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [5]),
        .Q(mscratch[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[6] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [6]),
        .Q(mscratch[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[7] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [7]),
        .Q(mscratch[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[8] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [8]),
        .Q(mscratch[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mscratch_reg[9] 
       (.C(clk),
        .CE(\mscratch[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [9]),
        .Q(mscratch[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[0] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [0]),
        .Q(mtime_compare[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[10] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [10]),
        .Q(mtime_compare[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[11] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [11]),
        .Q(mtime_compare[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[12] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [12]),
        .Q(mtime_compare[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[13] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [13]),
        .Q(mtime_compare[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[14] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [14]),
        .Q(mtime_compare[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[15] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [15]),
        .Q(mtime_compare[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[16] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [16]),
        .Q(mtime_compare[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[17] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [17]),
        .Q(mtime_compare[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[18] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [18]),
        .Q(mtime_compare[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[19] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [19]),
        .Q(mtime_compare[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[1] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [1]),
        .Q(mtime_compare[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[20] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [20]),
        .Q(mtime_compare[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[21] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [21]),
        .Q(mtime_compare[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[22] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [22]),
        .Q(mtime_compare[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[23] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [23]),
        .Q(mtime_compare[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[24] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [24]),
        .Q(mtime_compare[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[25] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [25]),
        .Q(mtime_compare[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[26] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [26]),
        .Q(mtime_compare[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[27] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [27]),
        .Q(mtime_compare[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[28] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [28]),
        .Q(mtime_compare[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[29] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [29]),
        .Q(mtime_compare[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[2] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [2]),
        .Q(mtime_compare[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[30] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [30]),
        .Q(mtime_compare[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[31] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [31]),
        .Q(mtime_compare[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[3] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [3]),
        .Q(mtime_compare[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[4] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [4]),
        .Q(mtime_compare[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[5] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [5]),
        .Q(mtime_compare[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[6] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [6]),
        .Q(mtime_compare[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[7] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [7]),
        .Q(mtime_compare[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[8] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [8]),
        .Q(mtime_compare[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtime_compare_reg[9] 
       (.C(clk),
        .CE(\mtime_compare[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [9]),
        .Q(mtime_compare[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(mtvec_out),
        .Q(\processor/mtvec [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[10]_i_1_n_0 ),
        .Q(\processor/mtvec [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[11]_i_1_n_0 ),
        .Q(\processor/mtvec [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[12]_i_1_n_0 ),
        .Q(\processor/mtvec [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[13]_i_1_n_0 ),
        .Q(\processor/mtvec [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[14]_i_1_n_0 ),
        .Q(\processor/mtvec [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[15]_i_1_n_0 ),
        .Q(\processor/mtvec [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[16]_i_1_n_0 ),
        .Q(\processor/mtvec [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[17]_i_1_n_0 ),
        .Q(\processor/mtvec [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[18]_i_1_n_0 ),
        .Q(\processor/mtvec [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[19]_i_1_n_0 ),
        .Q(\processor/mtvec [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[1]_i_1_n_0 ),
        .Q(\processor/mtvec [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[20]_i_1_n_0 ),
        .Q(\processor/mtvec [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[21]_i_1_n_0 ),
        .Q(\processor/mtvec [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[22]_i_1_n_0 ),
        .Q(\processor/mtvec [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[23]_i_1_n_0 ),
        .Q(\processor/mtvec [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[24]_i_1_n_0 ),
        .Q(\processor/mtvec [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[25]_i_1_n_0 ),
        .Q(\processor/mtvec [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[26]_i_1_n_0 ),
        .Q(\processor/mtvec [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[27]_i_1_n_0 ),
        .Q(\processor/mtvec [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[28]_i_1_n_0 ),
        .Q(\processor/mtvec [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[29]_i_1_n_0 ),
        .Q(\processor/mtvec [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[2]_i_1_n_0 ),
        .Q(\processor/mtvec [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[30]_i_1_n_0 ),
        .Q(\processor/mtvec [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[31]_i_1_n_0 ),
        .Q(\processor/mtvec [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[3]_i_1_n_0 ),
        .Q(\processor/mtvec [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[4]_i_1_n_0 ),
        .Q(\processor/mtvec [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[5]_i_1_n_0 ),
        .Q(\processor/mtvec [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[6]_i_1_n_0 ),
        .Q(\processor/mtvec [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[7]_i_1_n_0 ),
        .Q(\processor/mtvec [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[8]_i_1_n_0 ),
        .Q(\processor/mtvec [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_out_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\mtvec_out[9]_i_1_n_0 ),
        .Q(\processor/mtvec [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[0] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [0]),
        .Q(mtvec[0]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[10] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [10]),
        .Q(mtvec[10]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[11] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [11]),
        .Q(mtvec[11]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[12] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [12]),
        .Q(mtvec[12]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[13] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [13]),
        .Q(mtvec[13]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[14] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [14]),
        .Q(mtvec[14]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[15] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [15]),
        .Q(mtvec[15]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[16] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [16]),
        .Q(mtvec[16]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[17] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [17]),
        .Q(mtvec[17]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[18] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [18]),
        .Q(mtvec[18]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[19] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [19]),
        .Q(mtvec[19]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[1] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [1]),
        .Q(mtvec[1]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[20] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [20]),
        .Q(mtvec[20]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[21] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [21]),
        .Q(mtvec[21]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[22] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [22]),
        .Q(mtvec[22]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[23] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [23]),
        .Q(mtvec[23]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[24] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [24]),
        .Q(mtvec[24]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[25] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [25]),
        .Q(mtvec[25]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[26] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [26]),
        .Q(mtvec[26]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[27] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [27]),
        .Q(mtvec[27]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[28] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [28]),
        .Q(mtvec[28]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[29] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [29]),
        .Q(mtvec[29]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[2] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [2]),
        .Q(mtvec[2]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[30] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [30]),
        .Q(mtvec[30]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[31] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [31]),
        .Q(mtvec[31]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[3] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [3]),
        .Q(mtvec[3]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[4] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [4]),
        .Q(mtvec[4]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[5] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [5]),
        .Q(mtvec[5]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[6] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [6]),
        .Q(mtvec[6]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[7] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [7]),
        .Q(mtvec[7]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[8] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [8]),
        .Q(mtvec[8]),
        .S(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/mtvec_reg[9] 
       (.C(clk),
        .CE(\mtvec[31]_i_1_n_0 ),
        .D(\processor/wb_csr_data [9]),
        .Q(mtvec[9]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \processor/csr_unit/read_data_out2_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\processor/csr_unit/read_data_out2__3 ,\processor/csr_unit/read_data_out2_carry_n_1 ,\processor/csr_unit/read_data_out2_carry_n_2 ,\processor/csr_unit/read_data_out2_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({read_data_out2_carry_i_1_n_0,read_data_out2_carry_i_2_n_0,read_data_out2_carry_i_3_n_0,read_data_out2_carry_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(read_data_out),
        .Q(\processor/csr_read_data [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[10]_i_1_n_0 ),
        .Q(\processor/csr_read_data [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[11]_i_1_n_0 ),
        .Q(\processor/csr_read_data [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[12]_i_1_n_0 ),
        .Q(\processor/csr_read_data [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[13]_i_1_n_0 ),
        .Q(\processor/csr_read_data [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[14]_i_1_n_0 ),
        .Q(\processor/csr_read_data [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[15]_i_1_n_0 ),
        .Q(\processor/csr_read_data [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[16]_i_1_n_0 ),
        .Q(\processor/csr_read_data [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[17]_i_1_n_0 ),
        .Q(\processor/csr_read_data [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[18]_i_1_n_0 ),
        .Q(\processor/csr_read_data [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[19]_i_1_n_0 ),
        .Q(\processor/csr_read_data [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[1]_i_1_n_0 ),
        .Q(\processor/csr_read_data [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[20]_i_1_n_0 ),
        .Q(\processor/csr_read_data [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[21]_i_1_n_0 ),
        .Q(\processor/csr_read_data [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[22]_i_1_n_0 ),
        .Q(\processor/csr_read_data [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[23]_i_1_n_0 ),
        .Q(\processor/csr_read_data [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[24]_i_1_n_0 ),
        .Q(\processor/csr_read_data [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[25]_i_1_n_0 ),
        .Q(\processor/csr_read_data [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[26]_i_1_n_0 ),
        .Q(\processor/csr_read_data [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[27]_i_1_n_0 ),
        .Q(\processor/csr_read_data [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[28]_i_1_n_0 ),
        .Q(\processor/csr_read_data [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[29]_i_1_n_0 ),
        .Q(\processor/csr_read_data [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[2]_i_1_n_0 ),
        .Q(\processor/csr_read_data [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[30]_i_1_n_0 ),
        .Q(\processor/csr_read_data [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[31]_i_1_n_0 ),
        .Q(\processor/csr_read_data [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[3]_i_1_n_0 ),
        .Q(\processor/csr_read_data [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[4]_i_1_n_0 ),
        .Q(\processor/csr_read_data [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[5]_i_1_n_0 ),
        .Q(\processor/csr_read_data [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[6]_i_1_n_0 ),
        .Q(\processor/csr_read_data [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[7]_i_1_n_0 ),
        .Q(\processor/csr_read_data [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[8]_i_1_n_0 ),
        .Q(\processor/csr_read_data [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/read_data_out_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\read_data_out[9]_i_1_n_0 ),
        .Q(\processor/csr_read_data [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/software_interrupt_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(software_interrupt_i_1_n_0),
        .Q(\processor/software_interrupt ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[0] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[0]_i_1_n_7 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_ ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[10] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[8]_i_1_n_5 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[10] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[11] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[8]_i_1_n_4 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[11] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[12] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[12]_i_1_n_7 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[12] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[13] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[12]_i_1_n_6 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[13] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[14] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[12]_i_1_n_5 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[14] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[15] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[12]_i_1_n_4 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[15] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[16] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[16]_i_1_n_7 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[16] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[17] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[16]_i_1_n_6 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[17] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[18] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[16]_i_1_n_5 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[18] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[19] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[16]_i_1_n_4 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[19] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[1] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[0]_i_1_n_6 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[1] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[20] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[20]_i_1_n_7 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[20] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[21] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[20]_i_1_n_6 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[21] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[22] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[20]_i_1_n_5 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[22] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[23] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[20]_i_1_n_4 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[23] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[24] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[24]_i_1_n_7 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[24] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[25] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[24]_i_1_n_6 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[25] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[26] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[24]_i_1_n_5 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[26] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[27] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[24]_i_1_n_4 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[27] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[28] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[28]_i_1_n_7 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[28] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[29] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[28]_i_1_n_6 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[29] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[2] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[0]_i_1_n_5 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[2] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[30] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[28]_i_1_n_5 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[30] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[31] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[28]_i_1_n_4 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[31] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[32] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[32]_i_1_n_7 ),
        .Q(data12[0]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[33] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[32]_i_1_n_6 ),
        .Q(data12[1]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[34] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[32]_i_1_n_5 ),
        .Q(data12[2]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[35] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[32]_i_1_n_4 ),
        .Q(data12[3]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[36] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[36]_i_1_n_7 ),
        .Q(data12[4]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[37] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[36]_i_1_n_6 ),
        .Q(data12[5]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[38] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[36]_i_1_n_5 ),
        .Q(data12[6]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[39] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[36]_i_1_n_4 ),
        .Q(data12[7]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[3] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[0]_i_1_n_4 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[3] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[40] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[40]_i_1_n_7 ),
        .Q(data12[8]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[41] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[40]_i_1_n_6 ),
        .Q(data12[9]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[42] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[40]_i_1_n_5 ),
        .Q(data12[10]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[43] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[40]_i_1_n_4 ),
        .Q(data12[11]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[44] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[44]_i_1_n_7 ),
        .Q(data12[12]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[45] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[44]_i_1_n_6 ),
        .Q(data12[13]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[46] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[44]_i_1_n_5 ),
        .Q(data12[14]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[47] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[44]_i_1_n_4 ),
        .Q(data12[15]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[48] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[48]_i_1_n_7 ),
        .Q(data12[16]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[49] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[48]_i_1_n_6 ),
        .Q(data12[17]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[4] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[4]_i_1_n_7 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[4] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[50] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[48]_i_1_n_5 ),
        .Q(data12[18]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[51] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[48]_i_1_n_4 ),
        .Q(data12[19]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[52] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[52]_i_1_n_7 ),
        .Q(data12[20]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[53] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[52]_i_1_n_6 ),
        .Q(data12[21]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[54] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[52]_i_1_n_5 ),
        .Q(data12[22]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[55] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[52]_i_1_n_4 ),
        .Q(data12[23]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[56] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[56]_i_1_n_7 ),
        .Q(data12[24]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[57] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[56]_i_1_n_6 ),
        .Q(data12[25]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[58] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[56]_i_1_n_5 ),
        .Q(data12[26]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[59] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[56]_i_1_n_4 ),
        .Q(data12[27]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[5] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[4]_i_1_n_6 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[5] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[60] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[60]_i_1_n_7 ),
        .Q(data12[28]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[61] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[60]_i_1_n_6 ),
        .Q(data12[29]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[62] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[60]_i_1_n_5 ),
        .Q(data12[30]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[63] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[60]_i_1_n_4 ),
        .Q(data12[31]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[6] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[4]_i_1_n_5 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[6] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[7] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[4]_i_1_n_4 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[7] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[8] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[8]_i_1_n_7 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[8] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_counter/current_count_reg[9] 
       (.C(timer_clk),
        .CE(\<const1>__0__0 ),
        .D(\current_count_reg[8]_i_1_n_6 ),
        .Q(\processor/csr_unit/timer_counter/current_count_reg_n_0_[9] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \processor/csr_unit/timer_interrupt0_inferred__0_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\processor/csr_unit/timer_interrupt0_inferred__0_carry_n_0 ,\processor/csr_unit/timer_interrupt0_inferred__0_carry_n_1 ,\processor/csr_unit/timer_interrupt0_inferred__0_carry_n_2 ,\processor/csr_unit/timer_interrupt0_inferred__0_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({timer_interrupt0_inferred__0_carry_i_1_n_0,timer_interrupt0_inferred__0_carry_i_2_n_0,timer_interrupt0_inferred__0_carry_i_3_n_0,timer_interrupt0_inferred__0_carry_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \processor/csr_unit/timer_interrupt0_inferred__0_carry__0 
       (.CI(\processor/csr_unit/timer_interrupt0_inferred__0_carry_n_0 ),
        .CO({\processor/csr_unit/timer_interrupt0_inferred__0_carry__0_n_0 ,\processor/csr_unit/timer_interrupt0_inferred__0_carry__0_n_1 ,\processor/csr_unit/timer_interrupt0_inferred__0_carry__0_n_2 ,\processor/csr_unit/timer_interrupt0_inferred__0_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({timer_interrupt0_inferred__0_carry__0_i_1_n_0,timer_interrupt0_inferred__0_carry__0_i_2_n_0,timer_interrupt0_inferred__0_carry__0_i_3_n_0,timer_interrupt0_inferred__0_carry__0_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \processor/csr_unit/timer_interrupt0_inferred__0_carry__1 
       (.CI(\processor/csr_unit/timer_interrupt0_inferred__0_carry__0_n_0 ),
        .CO({\processor/csr_unit/timer_interrupt0_inferred__0_carry__1_n_0 ,\processor/csr_unit/timer_interrupt0_inferred__0_carry__1_n_1 ,\processor/csr_unit/timer_interrupt0_inferred__0_carry__1_n_2 ,\processor/csr_unit/timer_interrupt0_inferred__0_carry__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const0>__0__0 ,timer_interrupt0_inferred__0_carry__1_i_1_n_0,timer_interrupt0_inferred__0_carry__1_i_2_n_0,timer_interrupt0_inferred__0_carry__1_i_3_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/timer_interrupt_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(timer_interrupt_i_1_n_0),
        .Q(\processor/timer_interrupt ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[0] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [0]),
        .Q(tohost_data[0]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[10] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [10]),
        .Q(tohost_data[10]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[11] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [11]),
        .Q(tohost_data[11]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[12] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [12]),
        .Q(tohost_data[12]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[13] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [13]),
        .Q(tohost_data[13]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[14] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [14]),
        .Q(tohost_data[14]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[15] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [15]),
        .Q(tohost_data[15]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[16] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [16]),
        .Q(tohost_data[16]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[17] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [17]),
        .Q(tohost_data[17]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[18] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [18]),
        .Q(tohost_data[18]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[19] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [19]),
        .Q(tohost_data[19]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[1] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [1]),
        .Q(tohost_data[1]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[20] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [20]),
        .Q(tohost_data[20]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[21] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [21]),
        .Q(tohost_data[21]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[22] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [22]),
        .Q(tohost_data[22]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[23] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [23]),
        .Q(tohost_data[23]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[24] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [24]),
        .Q(tohost_data[24]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[25] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [25]),
        .Q(tohost_data[25]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[26] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [26]),
        .Q(tohost_data[26]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[27] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [27]),
        .Q(tohost_data[27]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[28] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [28]),
        .Q(tohost_data[28]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[29] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [29]),
        .Q(tohost_data[29]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[2] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [2]),
        .Q(tohost_data[2]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[30] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [30]),
        .Q(tohost_data[30]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[31] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [31]),
        .Q(tohost_data[31]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[3] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [3]),
        .Q(tohost_data[3]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[4] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [4]),
        .Q(tohost_data[4]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[5] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [5]),
        .Q(tohost_data[5]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[6] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [6]),
        .Q(tohost_data[6]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[7] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [7]),
        .Q(tohost_data[7]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[8] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [8]),
        .Q(tohost_data[8]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_data_reg[9] 
       (.C(clk),
        .CE(\processor/csr_unit/tohost_data0 ),
        .D(\processor/wb_csr_data [9]),
        .Q(tohost_data[9]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/csr_unit/tohost_updated_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\processor/csr_unit/tohost_data0 ),
        .Q(tohost_updated),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/count_instruction_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(count_instruction_i_1_n_0),
        .Q(\processor/id_count_instruction ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[10] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[10]),
        .Q(\processor/id_rd_address [3]),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[11] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[11]),
        .Q(\processor/id_rd_address [4]),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[12] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[12]),
        .Q(\processor/id_funct3 [0]),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[13] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[13]),
        .Q(\processor/id_funct3 [1]),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[14] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[14]),
        .Q(\processor/id_csr_use_immediate ),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[15] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[15]),
        .Q(\processor/id_rs1_address [0]),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[16] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[16]),
        .Q(\processor/id_rs1_address [1]),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[17] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[17]),
        .Q(\processor/id_rs1_address [2]),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[18] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[18]),
        .Q(\processor/id_rs1_address [3]),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[19] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[19]),
        .Q(\processor/id_rs1_address [4]),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[20] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[20]),
        .Q(\processor/id_shamt [0]),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[21] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[21]),
        .Q(\processor/id_shamt [1]),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[22] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[22]),
        .Q(\processor/id_shamt [2]),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[23] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[23]),
        .Q(\processor/id_shamt [3]),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[24] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[24]),
        .Q(\processor/id_shamt [4]),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[25] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[25]),
        .Q(data0[25]),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[26] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[26]),
        .Q(data0[26]),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[27] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[27]),
        .Q(data0[27]),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[28] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[28]),
        .Q(data0[28]),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[29] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[29]),
        .Q(data0[29]),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[2] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[2]),
        .Q(\processor/decode/instruction_reg_n_0_ ),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[30] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[30]),
        .Q(data0[30]),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[31] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[31]),
        .Q(data0[31]),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[3] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[3]),
        .Q(\processor/decode/instruction_reg_n_0_[3] ),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[4] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[4]),
        .Q(\processor/decode/instruction_reg_n_0_[4] ),
        .S(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[5] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[5]),
        .Q(\processor/decode/instruction_reg_n_0_[5] ),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[6] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[6]),
        .Q(\processor/decode/instruction_reg_n_0_[6] ),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[7] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[7]),
        .Q(\processor/id_rd_address [0]),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[8] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[8]),
        .Q(\processor/id_rd_address [1]),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/instruction_reg[9] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(imem_data[9]),
        .Q(\processor/id_rd_address [2]),
        .R(instruction));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[0] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[0]),
        .Q(\processor/id_pc [0]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[10] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[10]),
        .Q(\processor/id_pc [10]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[11] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[11]),
        .Q(\processor/id_pc [11]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[12] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[12]),
        .Q(\processor/id_pc [12]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[13] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[13]),
        .Q(\processor/id_pc [13]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[14] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[14]),
        .Q(\processor/id_pc [14]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[15] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[15]),
        .Q(\processor/id_pc [15]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[16] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[16]),
        .Q(\processor/id_pc [16]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[17] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[17]),
        .Q(\processor/id_pc [17]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[18] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[18]),
        .Q(\processor/id_pc [18]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[19] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[19]),
        .Q(\processor/id_pc [19]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[1] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[1]),
        .Q(\processor/id_pc [1]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[20] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[20]),
        .Q(\processor/id_pc [20]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[21] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[21]),
        .Q(\processor/id_pc [21]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[22] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[22]),
        .Q(\processor/id_pc [22]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[23] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[23]),
        .Q(\processor/id_pc [23]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[24] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[24]),
        .Q(\processor/id_pc [24]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[25] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[25]),
        .Q(\processor/id_pc [25]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[26] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[26]),
        .Q(\processor/id_pc [26]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[27] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[27]),
        .Q(\processor/id_pc [27]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[28] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[28]),
        .Q(\processor/id_pc [28]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[29] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[29]),
        .Q(\processor/id_pc [29]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[2] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[2]),
        .Q(\processor/id_pc [2]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[30] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[30]),
        .Q(\processor/id_pc [30]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[31] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[31]),
        .Q(\processor/id_pc [31]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[3] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[3]),
        .Q(\processor/id_pc [3]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[4] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[4]),
        .Q(\processor/id_pc [4]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[5] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[5]),
        .Q(\processor/id_pc [5]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[6] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[6]),
        .Q(\processor/id_pc [6]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[7] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[7]),
        .Q(\processor/id_pc [7]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/decode/pc_reg[8] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[8]),
        .Q(\processor/id_pc [8]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \processor/decode/pc_reg[9] 
       (.C(clk),
        .CE(\pc[31]_i_1_n_0 ),
        .D(pc[9]),
        .Q(\processor/id_pc [9]),
        .S(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[0] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [0]),
        .Q(dmem_address_p[0]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[10] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [10]),
        .Q(dmem_address_p[10]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[11] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [11]),
        .Q(dmem_address_p[11]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[12] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [12]),
        .Q(dmem_address_p[12]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[13] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [13]),
        .Q(dmem_address_p[13]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[14] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [14]),
        .Q(dmem_address_p[14]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[15] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [15]),
        .Q(dmem_address_p[15]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[16] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [16]),
        .Q(dmem_address_p[16]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[17] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [17]),
        .Q(dmem_address_p[17]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[18] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [18]),
        .Q(dmem_address_p[18]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[19] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [19]),
        .Q(dmem_address_p[19]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[1] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [1]),
        .Q(dmem_address_p[1]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[20] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [20]),
        .Q(dmem_address_p[20]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[21] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [21]),
        .Q(dmem_address_p[21]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[22] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [22]),
        .Q(dmem_address_p[22]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[23] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [23]),
        .Q(dmem_address_p[23]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[24] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [24]),
        .Q(dmem_address_p[24]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[25] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [25]),
        .Q(dmem_address_p[25]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[26] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [26]),
        .Q(dmem_address_p[26]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[27] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [27]),
        .Q(dmem_address_p[27]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[28] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [28]),
        .Q(dmem_address_p[28]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[29] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [29]),
        .Q(dmem_address_p[29]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[2] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [2]),
        .Q(dmem_address_p[2]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[30] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [30]),
        .Q(dmem_address_p[30]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[31] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [31]),
        .Q(dmem_address_p[31]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[3] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [3]),
        .Q(dmem_address_p[3]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[4] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [4]),
        .Q(dmem_address_p[4]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[5] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [5]),
        .Q(dmem_address_p[5]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[6] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [6]),
        .Q(dmem_address_p[6]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[7] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [7]),
        .Q(dmem_address_p[7]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[8] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [8]),
        .Q(dmem_address_p[8]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_address_p_reg[9] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_data [9]),
        .Q(dmem_address_p[9]),
        .R(\dmem_address_p[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[0] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [0]),
        .Q(dmem_data_out_p[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[10] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [10]),
        .Q(dmem_data_out_p[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[11] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [11]),
        .Q(dmem_data_out_p[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[12] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [12]),
        .Q(dmem_data_out_p[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[13] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [13]),
        .Q(dmem_data_out_p[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[14] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [14]),
        .Q(dmem_data_out_p[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[15] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [15]),
        .Q(dmem_data_out_p[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[16] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [16]),
        .Q(dmem_data_out_p[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[17] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [17]),
        .Q(dmem_data_out_p[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[18] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [18]),
        .Q(dmem_data_out_p[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[19] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [19]),
        .Q(dmem_data_out_p[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[1] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [1]),
        .Q(dmem_data_out_p[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[20] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [20]),
        .Q(dmem_data_out_p[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[21] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [21]),
        .Q(dmem_data_out_p[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[22] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [22]),
        .Q(dmem_data_out_p[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[23] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [23]),
        .Q(dmem_data_out_p[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[24] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [24]),
        .Q(dmem_data_out_p[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[25] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [25]),
        .Q(dmem_data_out_p[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[26] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [26]),
        .Q(dmem_data_out_p[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[27] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [27]),
        .Q(dmem_data_out_p[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[28] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [28]),
        .Q(dmem_data_out_p[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[29] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [29]),
        .Q(dmem_data_out_p[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[2] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [2]),
        .Q(dmem_data_out_p[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[30] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [30]),
        .Q(dmem_data_out_p[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[31] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [31]),
        .Q(dmem_data_out_p[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[3] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [3]),
        .Q(dmem_data_out_p[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[4] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [4]),
        .Q(dmem_data_out_p[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[5] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [5]),
        .Q(dmem_data_out_p[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[6] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [6]),
        .Q(dmem_data_out_p[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[7] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [7]),
        .Q(dmem_data_out_p[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[8] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [8]),
        .Q(dmem_data_out_p[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_out_p_reg[9] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_out [9]),
        .Q(dmem_data_out_p[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_size_p_reg[0] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_size [0]),
        .Q(\processor/dmem_data_size_p [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_data_size_p_reg[1] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_data_size [1]),
        .Q(\processor/dmem_data_size_p [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_read_req_p_reg 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_read_req ),
        .Q(\processor/dmem_read_req_p ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/dmem_write_req_p_reg 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_dmem_write_req ),
        .Q(\processor/dmem_write_req_p ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/alu_op_reg[0] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_alu_op [0]),
        .Q(\processor/execute/alu_op [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/alu_op_reg[1] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_alu_op [1]),
        .Q(\processor/execute/alu_op [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/alu_op_reg[2] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_alu_op [2]),
        .Q(\processor/execute/alu_op [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/alu_op_reg[3] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_alu_op [3]),
        .Q(\processor/execute/alu_op [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/alu_x_src_reg[0] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_alu_x_src [0]),
        .Q(\processor/execute/alu_x_src [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/alu_x_src_reg[1] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_alu_x_src [1]),
        .Q(\processor/execute/alu_x_src [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/alu_x_src_reg[2] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_alu_x_src [2]),
        .Q(\processor/execute/alu_x_src [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/alu_y_src_reg[0] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_alu_y_src [0]),
        .Q(\processor/execute/alu_y_src [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/alu_y_src_reg[1] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_alu_y_src [1]),
        .Q(\processor/execute/alu_y_src [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/alu_y_src_reg[2] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_alu_y_src [2]),
        .Q(\processor/execute/alu_y_src [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/branch_reg[0] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_branch [0]),
        .Q(\processor/ex_branch [0]),
        .R(\processor/execute/rd_write_out0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/branch_reg[1] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_branch [1]),
        .Q(\processor/ex_branch [1]),
        .R(\processor/execute/rd_write_out0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/branch_reg[2] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_branch [2]),
        .Q(\processor/ex_branch [2]),
        .R(\processor/execute/rd_write_out0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/count_instruction_out_reg 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_count_instruction ),
        .Q(\processor/ex_count_instruction ),
        .R(\processor/execute/rd_write_out0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/csr_addr_reg[0] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(csr_addr),
        .Q(\processor/ex_csr_address [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/csr_addr_reg[10] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\csr_addr[10]_i_1_n_0 ),
        .Q(\processor/ex_csr_address [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/csr_addr_reg[11] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\csr_addr[11]_i_1_n_0 ),
        .Q(\processor/ex_csr_address [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/csr_addr_reg[1] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\csr_addr[1]_i_1_n_0 ),
        .Q(\processor/ex_csr_address [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/csr_addr_reg[2] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\csr_addr[2]_i_1_n_0 ),
        .Q(\processor/ex_csr_address [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/csr_addr_reg[3] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\csr_addr[3]_i_1_n_0 ),
        .Q(\processor/ex_csr_address [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "processor/execute/csr_addr_reg[3]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/csr_addr_reg[3]_replica 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\csr_addr[3]_i_1_n_0 ),
        .Q(\processor/ex_csr_address[3]_repN ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/csr_addr_reg[4] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\csr_addr[4]_i_1_n_0 ),
        .Q(\processor/ex_csr_address [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/csr_addr_reg[5] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\csr_addr[5]_i_1_n_0 ),
        .Q(\processor/ex_csr_address [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/csr_addr_reg[6] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\csr_addr[6]_i_1_n_0 ),
        .Q(\processor/ex_csr_address [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "processor/execute/csr_addr_reg[6]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/csr_addr_reg[6]_replica 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\csr_addr[6]_i_1_n_0 ),
        .Q(\processor/ex_csr_address[6]_repN ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "processor/execute/csr_addr_reg[6]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/csr_addr_reg[6]_replica_1 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\csr_addr[6]_i_1_n_0 ),
        .Q(\processor/ex_csr_address[6]_repN_1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/csr_addr_reg[7] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\csr_addr[7]_i_1_n_0 ),
        .Q(\processor/ex_csr_address [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "processor/execute/csr_addr_reg[7]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/csr_addr_reg[7]_replica 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\csr_addr[7]_i_1_n_0 ),
        .Q(\processor/ex_csr_address[7]_repN ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/csr_addr_reg[8] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\csr_addr[8]_i_1_n_0 ),
        .Q(\processor/ex_csr_address [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/csr_addr_reg[9] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\csr_addr[9]_i_1_n_0 ),
        .Q(\processor/ex_csr_address [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/csr_write_reg[0] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_csr_write [0]),
        .Q(\processor/ex_csr_write [0]),
        .R(\processor/execute/rd_write_out0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/csr_write_reg[1] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_csr_write [1]),
        .Q(\processor/ex_csr_write [1]),
        .R(\processor/execute/rd_write_out0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/csr_writeable_reg 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/csr_read_writeable ),
        .Q(\processor/execute/csr_writeable ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/decode_exception_cause_reg[0] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_exception_cause [0]),
        .Q(\processor/execute/decode_exception_cause [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/decode_exception_cause_reg[2] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_exception_cause [2]),
        .Q(\processor/execute/decode_exception_cause [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/decode_exception_cause_reg[3] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_exception_cause [3]),
        .Q(\processor/execute/decode_exception_cause [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/decode_exception_reg 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_exception ),
        .Q(\processor/execute/decode_exception ),
        .R(\processor/execute/rd_write_out0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/funct3_reg[0] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_funct3 [0]),
        .Q(\processor/execute/funct3 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/funct3_reg[1] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_funct3 [1]),
        .Q(\processor/execute/funct3 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/funct3_reg[2] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_csr_use_immediate ),
        .Q(\processor/execute/funct3 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[0] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [0]),
        .Q(\processor/execute/immediate [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[10] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(data0[30]),
        .Q(\processor/execute/immediate [10]),
        .R(\immediate[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[11] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [11]),
        .Q(\processor/execute/immediate [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[12] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [12]),
        .Q(\processor/execute/immediate [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[13] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [13]),
        .Q(\processor/execute/immediate [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[14] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [14]),
        .Q(\processor/execute/immediate [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[15] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [15]),
        .Q(\processor/execute/immediate [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[16] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [16]),
        .Q(\processor/execute/immediate [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[17] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [17]),
        .Q(\processor/execute/immediate [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[18] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [18]),
        .Q(\processor/execute/immediate [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[19] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [19]),
        .Q(\processor/execute/immediate [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[1] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [1]),
        .Q(\processor/execute/immediate [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[20] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [20]),
        .Q(\processor/execute/immediate [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[21] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [21]),
        .Q(\processor/execute/immediate [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[22] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [22]),
        .Q(\processor/execute/immediate [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[23] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [23]),
        .Q(\processor/execute/immediate [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[24] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [24]),
        .Q(\processor/execute/immediate [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[25] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [25]),
        .Q(\processor/execute/immediate [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[26] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [26]),
        .Q(\processor/execute/immediate [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[27] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [27]),
        .Q(\processor/execute/immediate [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[28] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [28]),
        .Q(\processor/execute/immediate [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[29] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [29]),
        .Q(\processor/execute/immediate [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[2] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [2]),
        .Q(\processor/execute/immediate [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[30] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [30]),
        .Q(\processor/execute/immediate [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[31] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [31]),
        .Q(\processor/execute/immediate [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[3] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [3]),
        .Q(\processor/execute/immediate [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[4] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_immediate [4]),
        .Q(\processor/execute/immediate [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[5] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(data0[25]),
        .Q(\processor/execute/immediate [5]),
        .R(\immediate[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[6] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(data0[26]),
        .Q(\processor/execute/immediate [6]),
        .R(\immediate[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[7] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(data0[27]),
        .Q(\processor/execute/immediate [7]),
        .R(\immediate[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[8] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(data0[28]),
        .Q(\processor/execute/immediate [8]),
        .R(\immediate[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/immediate_reg[9] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(data0[29]),
        .Q(\processor/execute/immediate [9]),
        .R(\immediate[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mem_op_reg[0] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_mem_op [0]),
        .Q(\processor/ex_mem_op [0]),
        .R(\processor/execute/rd_write_out0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mem_op_reg[1] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\mem_op[1]_i_1_n_0 ),
        .Q(\processor/ex_mem_op [1]),
        .R(\processor/execute/rd_write_out0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mem_op_reg[2] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_mem_op [2]),
        .Q(\processor/ex_mem_op [2]),
        .R(\processor/execute/rd_write_out0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mem_size_reg[0] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_mem_size ),
        .Q(\processor/ex_dmem_data_size [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mem_size_reg[1] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\mem_size[1]_i_2_n_0 ),
        .Q(\processor/ex_mem_size ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mie_reg[24] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mie [24]),
        .Q(\processor/execute/mie [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mie_reg[25] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mie [25]),
        .Q(\processor/execute/mie [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mie_reg[26] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mie [26]),
        .Q(\processor/execute/mie [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mie_reg[27] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mie [27]),
        .Q(\processor/execute/mie [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mie_reg[28] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mie [28]),
        .Q(\processor/execute/mie [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mie_reg[29] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mie [29]),
        .Q(\processor/execute/mie [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mie_reg[30] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mie [30]),
        .Q(\processor/execute/mie [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mie_reg[31] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mie [31]),
        .Q(\processor/execute/mie [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mie_reg[3] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mie [3]),
        .Q(\processor/execute/mie [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mie_reg[7] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mie [7]),
        .Q(\processor/execute/mie [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[0] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [0]),
        .Q(\processor/execute/mtvec [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[10] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [10]),
        .Q(\processor/execute/mtvec [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[11] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [11]),
        .Q(\processor/execute/mtvec [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[12] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [12]),
        .Q(\processor/execute/mtvec [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[13] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [13]),
        .Q(\processor/execute/mtvec [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[14] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [14]),
        .Q(\processor/execute/mtvec [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[15] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [15]),
        .Q(\processor/execute/mtvec [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[16] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [16]),
        .Q(\processor/execute/mtvec [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[17] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [17]),
        .Q(\processor/execute/mtvec [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[18] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [18]),
        .Q(\processor/execute/mtvec [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[19] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [19]),
        .Q(\processor/execute/mtvec [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[1] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [1]),
        .Q(\processor/execute/mtvec [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[20] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [20]),
        .Q(\processor/execute/mtvec [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[21] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [21]),
        .Q(\processor/execute/mtvec [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[22] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [22]),
        .Q(\processor/execute/mtvec [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[23] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [23]),
        .Q(\processor/execute/mtvec [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[24] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [24]),
        .Q(\processor/execute/mtvec [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[25] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [25]),
        .Q(\processor/execute/mtvec [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[26] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [26]),
        .Q(\processor/execute/mtvec [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[27] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [27]),
        .Q(\processor/execute/mtvec [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[28] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [28]),
        .Q(\processor/execute/mtvec [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[29] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [29]),
        .Q(\processor/execute/mtvec [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[2] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [2]),
        .Q(\processor/execute/mtvec [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[30] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [30]),
        .Q(\processor/execute/mtvec [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[31] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [31]),
        .Q(\processor/execute/mtvec [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[3] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [3]),
        .Q(\processor/execute/mtvec [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[4] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [4]),
        .Q(\processor/execute/mtvec [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[5] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [5]),
        .Q(\processor/execute/mtvec [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[6] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [6]),
        .Q(\processor/execute/mtvec [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[7] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [7]),
        .Q(\processor/execute/mtvec [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[8] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [8]),
        .Q(\processor/execute/mtvec [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/mtvec_reg[9] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/mtvec [9]),
        .Q(\processor/execute/mtvec [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[0] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [0]),
        .Q(\processor/ex_pc [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[10] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [10]),
        .Q(\processor/ex_pc [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[11] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [11]),
        .Q(\processor/ex_pc [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[12] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [12]),
        .Q(\processor/ex_pc [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[13] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [13]),
        .Q(\processor/ex_pc [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[14] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [14]),
        .Q(\processor/ex_pc [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[15] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [15]),
        .Q(\processor/ex_pc [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[16] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [16]),
        .Q(\processor/ex_pc [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[17] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [17]),
        .Q(\processor/ex_pc [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[18] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [18]),
        .Q(\processor/ex_pc [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[19] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [19]),
        .Q(\processor/ex_pc [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[1] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [1]),
        .Q(\processor/ex_pc [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[20] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [20]),
        .Q(\processor/ex_pc [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[21] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [21]),
        .Q(\processor/ex_pc [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[22] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [22]),
        .Q(\processor/ex_pc [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[23] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [23]),
        .Q(\processor/ex_pc [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[24] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [24]),
        .Q(\processor/ex_pc [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[25] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [25]),
        .Q(\processor/ex_pc [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[26] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [26]),
        .Q(\processor/ex_pc [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[27] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [27]),
        .Q(\processor/ex_pc [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[28] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [28]),
        .Q(\processor/ex_pc [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[29] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [29]),
        .Q(\processor/ex_pc [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[2] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [2]),
        .Q(\processor/ex_pc [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[30] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [30]),
        .Q(\processor/ex_pc [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[31] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [31]),
        .Q(\processor/ex_pc [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[3] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [3]),
        .Q(\processor/ex_pc [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[4] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [4]),
        .Q(\processor/ex_pc [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[5] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [5]),
        .Q(\processor/ex_pc [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[6] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [6]),
        .Q(\processor/ex_pc [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[7] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [7]),
        .Q(\processor/ex_pc [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[8] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [8]),
        .Q(\processor/ex_pc [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/pc_reg[9] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_pc [9]),
        .Q(\processor/ex_pc [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/rd_addr_out_reg[0] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_rd_address [0]),
        .Q(\processor/ex_rd_address [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/rd_addr_out_reg[1] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_rd_address [1]),
        .Q(\processor/ex_rd_address [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/rd_addr_out_reg[2] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_rd_address [2]),
        .Q(\processor/ex_rd_address [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/rd_addr_out_reg[3] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_rd_address [3]),
        .Q(\processor/ex_rd_address [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/rd_addr_out_reg[4] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_rd_address [4]),
        .Q(\processor/ex_rd_address [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/rd_write_out_reg 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_rd_write ),
        .Q(\processor/ex_rd_write ),
        .R(\processor/execute/rd_write_out0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/rs1_addr_reg[0] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/rs1_address [0]),
        .Q(\processor/execute/rs1_addr [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "processor/execute/rs1_addr_reg[0]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/rs1_addr_reg[0]_replica 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/rs1_address [0]),
        .Q(\processor/execute/rs1_addr[0]_repN ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/rs1_addr_reg[1] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/rs1_address [1]),
        .Q(\processor/execute/rs1_addr [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/rs1_addr_reg[2] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/rs1_address [2]),
        .Q(\processor/execute/rs1_addr [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/rs1_addr_reg[3] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/rs1_address [3]),
        .Q(\processor/execute/rs1_addr [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/rs1_addr_reg[4] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/rs1_address [4]),
        .Q(\processor/execute/rs1_addr [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/rs2_addr_reg[0] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/rs2_address [0]),
        .Q(\processor/execute/rs2_addr [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/rs2_addr_reg[1] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/rs2_address [1]),
        .Q(\processor/execute/rs2_addr [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/rs2_addr_reg[2] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/rs2_address [2]),
        .Q(\processor/execute/rs2_addr [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/rs2_addr_reg[3] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/rs2_address [3]),
        .Q(\processor/execute/rs2_addr [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/rs2_addr_reg[4] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/rs2_address [4]),
        .Q(\processor/execute/rs2_addr [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/shamt_reg[0] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_shamt [0]),
        .Q(\processor/execute/shamt [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/shamt_reg[1] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_shamt [1]),
        .Q(\processor/execute/shamt [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/shamt_reg[2] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_shamt [2]),
        .Q(\processor/execute/shamt [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/shamt_reg[3] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_shamt [3]),
        .Q(\processor/execute/shamt [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/execute/shamt_reg[4] 
       (.C(clk),
        .CE(\mem_size[1]_i_1_n_0 ),
        .D(\processor/id_shamt [4]),
        .Q(\processor/execute/shamt [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/cancel_fetch_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(cancel_fetch_i_1_n_0),
        .Q(\processor/fetch/cancel_fetch ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[0] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[0]),
        .Q(pc[0]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[10] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[10]),
        .Q(pc[10]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[11] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[11]),
        .Q(pc[11]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[12] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[12]),
        .Q(pc[12]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[13] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[13]),
        .Q(pc[13]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[14] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[14]),
        .Q(pc[14]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[15] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[15]),
        .Q(pc[15]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[16] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[16]),
        .Q(pc[16]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[17] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[17]),
        .Q(pc[17]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[18] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[18]),
        .Q(pc[18]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[19] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[19]),
        .Q(pc[19]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[1] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[1]),
        .Q(pc[1]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[20] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[20]),
        .Q(pc[20]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[21] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[21]),
        .Q(pc[21]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[22] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[22]),
        .Q(pc[22]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[23] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[23]),
        .Q(pc[23]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[24] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[24]),
        .Q(pc[24]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[25] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[25]),
        .Q(pc[25]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[26] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[26]),
        .Q(pc[26]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[27] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[27]),
        .Q(pc[27]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[28] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[28]),
        .Q(pc[28]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[29] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[29]),
        .Q(pc[29]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[2] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[2]),
        .Q(pc[2]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[30] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[30]),
        .Q(pc[30]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[31] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[31]),
        .Q(pc[31]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[3] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[3]),
        .Q(pc[3]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[4] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[4]),
        .Q(pc[4]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[5] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[5]),
        .Q(pc[5]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[6] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[6]),
        .Q(pc[6]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[7] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[7]),
        .Q(pc[7]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[8] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[8]),
        .Q(pc[8]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \processor/fetch/pc_reg[9] 
       (.C(clk),
        .CE(\pc[31]_i_1__0_n_0 ),
        .D(pc_next[9]),
        .Q(pc[9]),
        .S(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/count_instr_out_reg 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_count_instruction ),
        .Q(count_instr_out),
        .R(count_instr_out_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \processor/memory/csr_addr_out_reg[0] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_csr_address [0]),
        .Q(\processor/mem_csr_address [0]),
        .S(csr_addr_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_addr_out_reg[10] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_csr_address [10]),
        .Q(\processor/mem_csr_address [10]),
        .R(csr_addr_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_addr_out_reg[11] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_csr_address [11]),
        .Q(\processor/mem_csr_address [11]),
        .R(csr_addr_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_addr_out_reg[1] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_csr_address [1]),
        .Q(\processor/mem_csr_address [1]),
        .R(csr_addr_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_addr_out_reg[2] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_csr_address [2]),
        .Q(\processor/mem_csr_address [2]),
        .R(csr_addr_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_addr_out_reg[3] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_csr_address [3]),
        .Q(\processor/mem_csr_address [3]),
        .R(csr_addr_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_addr_out_reg[4] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_csr_address [4]),
        .Q(\processor/mem_csr_address [4]),
        .R(csr_addr_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "processor/memory/csr_addr_out_reg[4]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_addr_out_reg[4]_replica 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_csr_address [4]),
        .Q(\processor/mem_csr_address[4]_repN ),
        .R(csr_addr_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "processor/memory/csr_addr_out_reg[4]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_addr_out_reg[4]_replica_1 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_csr_address [4]),
        .Q(\processor/mem_csr_address[4]_repN_1 ),
        .R(csr_addr_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_addr_out_reg[5] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_csr_address [5]),
        .Q(\processor/mem_csr_address [5]),
        .R(csr_addr_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \processor/memory/csr_addr_out_reg[6] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_csr_address [6]),
        .Q(\processor/mem_csr_address [6]),
        .S(csr_addr_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_addr_out_reg[7] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_csr_address [7]),
        .Q(\processor/mem_csr_address [7]),
        .R(csr_addr_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \processor/memory/csr_addr_out_reg[8] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_csr_address [8]),
        .Q(\processor/mem_csr_address [8]),
        .S(csr_addr_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \processor/memory/csr_addr_out_reg[9] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_csr_address [9]),
        .Q(\processor/mem_csr_address [9]),
        .S(csr_addr_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[0] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(csr_data_out),
        .Q(\processor/mem_csr_data [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[10] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[10]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[11] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[11]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[12] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[12]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[13] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[13]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[14] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[14]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[15] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[15]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[16] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[16]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[17] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[17]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[18] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[18]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[19] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[19]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[1] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[1]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[20] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[20]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[21] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[21]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[22] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[22]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[23] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[23]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[24] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[24]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[25] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[25]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[26] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[26]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[27] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[27]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[28] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[28]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[29] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[29]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[2] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[2]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[30] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[30]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[31] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[31]_i_2_n_0 ),
        .Q(\processor/mem_csr_data [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[3] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[3]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[4] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[4]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[5] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[5]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[6] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[6]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[7] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[7]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[8] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[8]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_data_out_reg[9] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\csr_data_out[9]_i_1_n_0 ),
        .Q(\processor/mem_csr_data [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEFE0)) 
    \processor/memory/csr_write_out[0]_i_1 
       (.I0(\processor/ex_csr_write [0]),
        .I1(\mem_op[2]_i_5_n_0 ),
        .I2(\processor/memory/p_1_in ),
        .I3(\processor/mem_csr_write [0]),
        .O(\processor/memory/csr_write_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEFE0)) 
    \processor/memory/csr_write_out[1]_i_1 
       (.I0(\processor/ex_csr_write [1]),
        .I1(\mem_op[2]_i_5_n_0 ),
        .I2(\processor/memory/p_1_in ),
        .I3(\processor/mem_csr_write [1]),
        .O(\processor/memory/csr_write_out[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_write_out_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\processor/memory/csr_write_out ),
        .Q(\processor/mem_csr_write [0]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/csr_write_out_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\processor/memory/csr_write_out[1]_i_1_n_0 ),
        .Q(\processor/mem_csr_write [1]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][0] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [0]),
        .Q(\processor/mem_exception_context[badaddr] [0]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][10] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [10]),
        .Q(\processor/mem_exception_context[badaddr] [10]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][11] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [11]),
        .Q(\processor/mem_exception_context[badaddr] [11]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][12] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [12]),
        .Q(\processor/mem_exception_context[badaddr] [12]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][13] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [13]),
        .Q(\processor/mem_exception_context[badaddr] [13]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][14] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [14]),
        .Q(\processor/mem_exception_context[badaddr] [14]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][15] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [15]),
        .Q(\processor/mem_exception_context[badaddr] [15]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][16] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [16]),
        .Q(\processor/mem_exception_context[badaddr] [16]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][17] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [17]),
        .Q(\processor/mem_exception_context[badaddr] [17]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][18] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [18]),
        .Q(\processor/mem_exception_context[badaddr] [18]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][19] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [19]),
        .Q(\processor/mem_exception_context[badaddr] [19]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][1] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [1]),
        .Q(\processor/mem_exception_context[badaddr] [1]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][20] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [20]),
        .Q(\processor/mem_exception_context[badaddr] [20]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][21] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [21]),
        .Q(\processor/mem_exception_context[badaddr] [21]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][22] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [22]),
        .Q(\processor/mem_exception_context[badaddr] [22]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][23] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [23]),
        .Q(\processor/mem_exception_context[badaddr] [23]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][24] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [24]),
        .Q(\processor/mem_exception_context[badaddr] [24]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][25] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [25]),
        .Q(\processor/mem_exception_context[badaddr] [25]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][26] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [26]),
        .Q(\processor/mem_exception_context[badaddr] [26]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][27] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [27]),
        .Q(\processor/mem_exception_context[badaddr] [27]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][28] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [28]),
        .Q(\processor/mem_exception_context[badaddr] [28]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][29] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [29]),
        .Q(\processor/mem_exception_context[badaddr] [29]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][2] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [2]),
        .Q(\processor/mem_exception_context[badaddr] [2]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][30] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [30]),
        .Q(\processor/mem_exception_context[badaddr] [30]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][31] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [31]),
        .Q(\processor/mem_exception_context[badaddr] [31]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][3] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [3]),
        .Q(\processor/mem_exception_context[badaddr] [3]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][4] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [4]),
        .Q(\processor/mem_exception_context[badaddr] [4]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][5] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [5]),
        .Q(\processor/mem_exception_context[badaddr] [5]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][6] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [6]),
        .Q(\processor/mem_exception_context[badaddr] [6]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][7] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [7]),
        .Q(\processor/mem_exception_context[badaddr] [7]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][8] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [8]),
        .Q(\processor/mem_exception_context[badaddr] [8]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[badaddr][9] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[badaddr] [9]),
        .Q(\processor/mem_exception_context[badaddr] [9]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[cause][0] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[cause] [0]),
        .Q(\processor/mem_exception_context[cause] [0]),
        .S(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[cause][1] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[cause] [1]),
        .Q(\processor/mem_exception_context[cause] [1]),
        .S(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[cause][2] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[cause] [2]),
        .Q(\processor/mem_exception_context[cause] [2]),
        .S(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[cause][3] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[cause] [3]),
        .Q(\processor/mem_exception_context[cause] [3]),
        .S(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[cause][4] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[cause] [4]),
        .Q(\processor/mem_exception_context[cause] [4]),
        .S(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[cause][5] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/ex_exception_context[cause] [5]),
        .Q(\processor/mem_exception_context[cause] [5]),
        .R(\exception_context_out[badaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[ie1] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\exception_context_out[ie1]_i_1_n_0 ),
        .Q(\processor/mem_exception_context ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_context_out_reg[ie] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\exception_context_out[ie]_i_1_n_0 ),
        .Q(\processor/mem_exception_context[ie] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/exception_out_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\processor/memory/exception_out0 ),
        .Q(\processor/mem_exception ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/mem_op_reg[0] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_mem_op [0]),
        .Q(\processor/mem_mem_op [0]),
        .R(count_instr_out_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/mem_op_reg[1] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_mem_op [1]),
        .Q(\processor/mem_mem_op [1]),
        .R(count_instr_out_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "processor/memory/mem_op_reg[1]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/mem_op_reg[1]_replica 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_mem_op [1]),
        .Q(\processor/mem_mem_op[1]_repN ),
        .R(count_instr_out_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "processor/memory/mem_op_reg[1]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/mem_op_reg[1]_replica_1 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_mem_op [1]),
        .Q(\processor/mem_mem_op[1]_repN_1 ),
        .R(count_instr_out_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "processor/memory/mem_op_reg[1]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/mem_op_reg[1]_replica_2 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_mem_op [1]),
        .Q(\processor/mem_mem_op[1]_repN_2 ),
        .R(count_instr_out_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/mem_op_reg[2] 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_mem_op [2]),
        .Q(\processor/mem_mem_op [2]),
        .R(count_instr_out_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/mem_size_reg[0] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_dmem_data_size [1]),
        .Q(mem_size[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "processor/memory/mem_size_reg[0]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/mem_size_reg[0]_replica 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_dmem_data_size [1]),
        .Q(\mem_size[0]_repN ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/mem_size_reg[1] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_mem_size ),
        .Q(mem_size[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "processor/memory/mem_size_reg[1]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/mem_size_reg[1]_replica 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_mem_size ),
        .Q(\mem_size[1]_repN ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "processor/memory/mem_size_reg[1]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/mem_size_reg[1]_replica_1 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_mem_size ),
        .Q(\mem_size[1]_repN_1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "processor/memory/mem_size_reg[1]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/mem_size_reg[1]_replica_2 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_mem_size ),
        .Q(\mem_size[1]_repN_2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_addr_out_reg[0] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_address [0]),
        .Q(\processor/mem_rd_address [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_addr_out_reg[1] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_address [1]),
        .Q(\processor/mem_rd_address [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_addr_out_reg[2] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_address [2]),
        .Q(\processor/mem_rd_address [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_addr_out_reg[3] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_address [3]),
        .Q(\processor/mem_rd_address [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_addr_out_reg[4] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_address [4]),
        .Q(\processor/mem_rd_address [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[0] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [0]),
        .Q(rd_data[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[10] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [10]),
        .Q(rd_data[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[11] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [11]),
        .Q(rd_data[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[12] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [12]),
        .Q(rd_data[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[13] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [13]),
        .Q(rd_data[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[14] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [14]),
        .Q(rd_data[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[15] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [15]),
        .Q(rd_data[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[16] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [16]),
        .Q(rd_data[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[17] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [17]),
        .Q(rd_data[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[18] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [18]),
        .Q(rd_data[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[19] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [19]),
        .Q(rd_data[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[1] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [1]),
        .Q(rd_data[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[20] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [20]),
        .Q(rd_data[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[21] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [21]),
        .Q(rd_data[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[22] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [22]),
        .Q(rd_data[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[23] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [23]),
        .Q(rd_data[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[24] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [24]),
        .Q(rd_data[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[25] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [25]),
        .Q(rd_data[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[26] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [26]),
        .Q(rd_data[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[27] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [27]),
        .Q(rd_data[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[28] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [28]),
        .Q(rd_data[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[29] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [29]),
        .Q(rd_data[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[2] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [2]),
        .Q(rd_data[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[30] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [30]),
        .Q(rd_data[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[31] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [31]),
        .Q(rd_data[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[3] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [3]),
        .Q(rd_data[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[4] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [4]),
        .Q(rd_data[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[5] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [5]),
        .Q(rd_data[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[6] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [6]),
        .Q(rd_data[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[7] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [7]),
        .Q(rd_data[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[8] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [8]),
        .Q(rd_data[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_data_reg[9] 
       (.C(clk),
        .CE(\csr_data_out[31]_i_1_n_0 ),
        .D(\processor/ex_rd_data [9]),
        .Q(rd_data[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/memory/rd_write_out_reg 
       (.C(clk),
        .CE(\processor/memory/p_1_in ),
        .D(\processor/ex_rd_write ),
        .Q(\processor/mem_rd_write ),
        .R(count_instr_out_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \processor/regfile/registers_reg_r1_0_31_0_5 
       (.ADDRA(\processor/rs2_address ),
        .ADDRB(\processor/rs2_address ),
        .ADDRC(\processor/rs2_address ),
        .ADDRD(\processor/wb_rd_address ),
        .DIA(\processor/wb_rd_data [1:0]),
        .DIB(\processor/wb_rd_data [3:2]),
        .DIC(\processor/wb_rd_data [5:4]),
        .DID({\<const0>__0__0 ,\<const0>__0__0 }),
        .DOA(p_2_out[1:0]),
        .DOB(p_2_out[3:2]),
        .DOC(p_2_out[5:4]),
        .WCLK(clk),
        .WE(\processor/regfile/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \processor/regfile/registers_reg_r1_0_31_12_17 
       (.ADDRA(\processor/rs2_address ),
        .ADDRB(\processor/rs2_address ),
        .ADDRC(\processor/rs2_address ),
        .ADDRD(\processor/wb_rd_address ),
        .DIA(\processor/wb_rd_data [13:12]),
        .DIB(\processor/wb_rd_data [15:14]),
        .DIC(\processor/wb_rd_data [17:16]),
        .DID({\<const0>__0__0 ,\<const0>__0__0 }),
        .DOA(p_2_out[13:12]),
        .DOB(p_2_out[15:14]),
        .DOC(p_2_out[17:16]),
        .WCLK(clk),
        .WE(\processor/regfile/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \processor/regfile/registers_reg_r1_0_31_18_23 
       (.ADDRA(\processor/rs2_address ),
        .ADDRB(\processor/rs2_address ),
        .ADDRC(\processor/rs2_address ),
        .ADDRD(\processor/wb_rd_address ),
        .DIA(\processor/wb_rd_data [19:18]),
        .DIB(\processor/wb_rd_data [21:20]),
        .DIC(\processor/wb_rd_data [23:22]),
        .DID({\<const0>__0__0 ,\<const0>__0__0 }),
        .DOA(p_2_out[19:18]),
        .DOB(p_2_out[21:20]),
        .DOC(p_2_out[23:22]),
        .WCLK(clk),
        .WE(\processor/regfile/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \processor/regfile/registers_reg_r1_0_31_24_29 
       (.ADDRA(\processor/rs2_address ),
        .ADDRB(\processor/rs2_address ),
        .ADDRC(\processor/rs2_address ),
        .ADDRD(\processor/wb_rd_address ),
        .DIA(\processor/wb_rd_data [25:24]),
        .DIB(\processor/wb_rd_data [27:26]),
        .DIC(\processor/wb_rd_data [29:28]),
        .DID({\<const0>__0__0 ,\<const0>__0__0 }),
        .DOA(p_2_out[25:24]),
        .DOB(p_2_out[27:26]),
        .DOC(p_2_out[29:28]),
        .WCLK(clk),
        .WE(\processor/regfile/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \processor/regfile/registers_reg_r1_0_31_30_31 
       (.ADDRA(\processor/rs2_address ),
        .ADDRB(\processor/rs2_address ),
        .ADDRC(\processor/rs2_address ),
        .ADDRD(\processor/wb_rd_address ),
        .DIA(\processor/wb_rd_data [31:30]),
        .DIB({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIC({\<const0>__0__0 ,\<const0>__0__0 }),
        .DID({\<const0>__0__0 ,\<const0>__0__0 }),
        .DOA(p_2_out[31:30]),
        .WCLK(clk),
        .WE(\processor/regfile/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \processor/regfile/registers_reg_r1_0_31_6_11 
       (.ADDRA(\processor/rs2_address ),
        .ADDRB(\processor/rs2_address ),
        .ADDRC(\processor/rs2_address ),
        .ADDRD(\processor/wb_rd_address ),
        .DIA(\processor/wb_rd_data [7:6]),
        .DIB(\processor/wb_rd_data [9:8]),
        .DIC(\processor/wb_rd_data [11:10]),
        .DID({\<const0>__0__0 ,\<const0>__0__0 }),
        .DOA(p_2_out[7:6]),
        .DOB(p_2_out[9:8]),
        .DOC(p_2_out[11:10]),
        .WCLK(clk),
        .WE(\processor/regfile/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \processor/regfile/registers_reg_r2_0_31_0_5 
       (.ADDRA(\processor/rs1_address ),
        .ADDRB(\processor/rs1_address ),
        .ADDRC(\processor/rs1_address ),
        .ADDRD(\processor/wb_rd_address ),
        .DIA(\processor/wb_rd_data [1:0]),
        .DIB(\processor/wb_rd_data [3:2]),
        .DIC(\processor/wb_rd_data [5:4]),
        .DID({\<const0>__0__0 ,\<const0>__0__0 }),
        .DOA(p_1_out0_in[1:0]),
        .DOB(p_1_out0_in[3:2]),
        .DOC(p_1_out0_in[5:4]),
        .WCLK(clk),
        .WE(\processor/regfile/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \processor/regfile/registers_reg_r2_0_31_12_17 
       (.ADDRA(\processor/rs1_address ),
        .ADDRB(\processor/rs1_address ),
        .ADDRC(\processor/rs1_address ),
        .ADDRD(\processor/wb_rd_address ),
        .DIA(\processor/wb_rd_data [13:12]),
        .DIB(\processor/wb_rd_data [15:14]),
        .DIC(\processor/wb_rd_data [17:16]),
        .DID({\<const0>__0__0 ,\<const0>__0__0 }),
        .DOA(p_1_out0_in[13:12]),
        .DOB(p_1_out0_in[15:14]),
        .DOC(p_1_out0_in[17:16]),
        .WCLK(clk),
        .WE(\processor/regfile/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \processor/regfile/registers_reg_r2_0_31_18_23 
       (.ADDRA(\processor/rs1_address ),
        .ADDRB(\processor/rs1_address ),
        .ADDRC(\processor/rs1_address ),
        .ADDRD(\processor/wb_rd_address ),
        .DIA(\processor/wb_rd_data [19:18]),
        .DIB(\processor/wb_rd_data [21:20]),
        .DIC(\processor/wb_rd_data [23:22]),
        .DID({\<const0>__0__0 ,\<const0>__0__0 }),
        .DOA(p_1_out0_in[19:18]),
        .DOB(p_1_out0_in[21:20]),
        .DOC(p_1_out0_in[23:22]),
        .WCLK(clk),
        .WE(\processor/regfile/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \processor/regfile/registers_reg_r2_0_31_24_29 
       (.ADDRA(\processor/rs1_address ),
        .ADDRB(\processor/rs1_address ),
        .ADDRC(\processor/rs1_address ),
        .ADDRD(\processor/wb_rd_address ),
        .DIA(\processor/wb_rd_data [25:24]),
        .DIB(\processor/wb_rd_data [27:26]),
        .DIC(\processor/wb_rd_data [29:28]),
        .DID({\<const0>__0__0 ,\<const0>__0__0 }),
        .DOA(p_1_out0_in[25:24]),
        .DOB(p_1_out0_in[27:26]),
        .DOC(p_1_out0_in[29:28]),
        .WCLK(clk),
        .WE(\processor/regfile/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \processor/regfile/registers_reg_r2_0_31_30_31 
       (.ADDRA(\processor/rs1_address ),
        .ADDRB(\processor/rs1_address ),
        .ADDRC(\processor/rs1_address ),
        .ADDRD(\processor/wb_rd_address ),
        .DIA(\processor/wb_rd_data [31:30]),
        .DIB({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIC({\<const0>__0__0 ,\<const0>__0__0 }),
        .DID({\<const0>__0__0 ,\<const0>__0__0 }),
        .DOA(p_1_out0_in[31:30]),
        .WCLK(clk),
        .WE(\processor/regfile/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \processor/regfile/registers_reg_r2_0_31_6_11 
       (.ADDRA(\processor/rs1_address ),
        .ADDRB(\processor/rs1_address ),
        .ADDRC(\processor/rs1_address ),
        .ADDRD(\processor/wb_rd_address ),
        .DIA(\processor/wb_rd_data [7:6]),
        .DIB(\processor/wb_rd_data [9:8]),
        .DIC(\processor/wb_rd_data [11:10]),
        .DID({\<const0>__0__0 ,\<const0>__0__0 }),
        .DOA(p_1_out0_in[7:6]),
        .DOB(p_1_out0_in[9:8]),
        .DOC(p_1_out0_in[11:10]),
        .WCLK(clk),
        .WE(\processor/regfile/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[0]),
        .Q(\processor/rs1_data [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[10]),
        .Q(\processor/rs1_data [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[11]),
        .Q(\processor/rs1_data [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[12]),
        .Q(\processor/rs1_data [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[13]),
        .Q(\processor/rs1_data [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[14]),
        .Q(\processor/rs1_data [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[15]),
        .Q(\processor/rs1_data [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[16]),
        .Q(\processor/rs1_data [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[17]),
        .Q(\processor/rs1_data [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[18]),
        .Q(\processor/rs1_data [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[19]),
        .Q(\processor/rs1_data [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[1]),
        .Q(\processor/rs1_data [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[20]),
        .Q(\processor/rs1_data [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[21]),
        .Q(\processor/rs1_data [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[22]),
        .Q(\processor/rs1_data [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[23]),
        .Q(\processor/rs1_data [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[24]),
        .Q(\processor/rs1_data [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[25]),
        .Q(\processor/rs1_data [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[26]),
        .Q(\processor/rs1_data [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[27]),
        .Q(\processor/rs1_data [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[28]),
        .Q(\processor/rs1_data [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[29]),
        .Q(\processor/rs1_data [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[2]),
        .Q(\processor/rs1_data [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[30]),
        .Q(\processor/rs1_data [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[31]),
        .Q(\processor/rs1_data [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[3]),
        .Q(\processor/rs1_data [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[4]),
        .Q(\processor/rs1_data [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[5]),
        .Q(\processor/rs1_data [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[6]),
        .Q(\processor/rs1_data [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[7]),
        .Q(\processor/rs1_data [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[8]),
        .Q(\processor/rs1_data [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs1_data_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_1_out2_out[9]),
        .Q(\processor/rs1_data [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[0]),
        .Q(\processor/rs2_data [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[10]),
        .Q(\processor/rs2_data [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[11]),
        .Q(\processor/rs2_data [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[12]),
        .Q(\processor/rs2_data [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[13]),
        .Q(\processor/rs2_data [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[14]),
        .Q(\processor/rs2_data [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[15]),
        .Q(\processor/rs2_data [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[16]),
        .Q(\processor/rs2_data [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[17]),
        .Q(\processor/rs2_data [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[18]),
        .Q(\processor/rs2_data [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[19]),
        .Q(\processor/rs2_data [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[1]),
        .Q(\processor/rs2_data [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[20]),
        .Q(\processor/rs2_data [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[21]),
        .Q(\processor/rs2_data [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[22]),
        .Q(\processor/rs2_data [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[23]),
        .Q(\processor/rs2_data [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[24]),
        .Q(\processor/rs2_data [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[25]),
        .Q(\processor/rs2_data [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[26]),
        .Q(\processor/rs2_data [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[27]),
        .Q(\processor/rs2_data [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[28]),
        .Q(\processor/rs2_data [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[29]),
        .Q(\processor/rs2_data [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[2]),
        .Q(\processor/rs2_data [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[30]),
        .Q(\processor/rs2_data [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[31]),
        .Q(\processor/rs2_data [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[3]),
        .Q(\processor/rs2_data [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[4]),
        .Q(\processor/rs2_data [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[5]),
        .Q(\processor/rs2_data [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[6]),
        .Q(\processor/rs2_data [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[7]),
        .Q(\processor/rs2_data [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[8]),
        .Q(\processor/rs2_data [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/regfile/rs2_data_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_0_out1_out[9]),
        .Q(\processor/rs2_data [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/rs1_address_p_reg[0] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_rs1_address [0]),
        .Q(\processor/rs1_address_p [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/rs1_address_p_reg[1] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_rs1_address [1]),
        .Q(\processor/rs1_address_p [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/rs1_address_p_reg[2] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_rs1_address [2]),
        .Q(\processor/rs1_address_p [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/rs1_address_p_reg[3] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_rs1_address [3]),
        .Q(\processor/rs1_address_p [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/rs1_address_p_reg[4] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_rs1_address [4]),
        .Q(\processor/rs1_address_p [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/rs2_address_p_reg[0] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_shamt [0]),
        .Q(\processor/rs2_address_p [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/rs2_address_p_reg[1] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_shamt [1]),
        .Q(\processor/rs2_address_p [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/rs2_address_p_reg[2] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_shamt [2]),
        .Q(\processor/rs2_address_p [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/rs2_address_p_reg[3] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_shamt [3]),
        .Q(\processor/rs2_address_p [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/rs2_address_p_reg[4] 
       (.C(clk),
        .CE(\processor/execute/exception_taken0 ),
        .D(\processor/id_shamt [4]),
        .Q(\processor/rs2_address_p [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/count_instr_out_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(count_instr_out),
        .Q(\processor/writeback/count_instr_out_reg_n_0 ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_addr_out_reg[0] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_address [0]),
        .Q(\processor/wb_csr_address [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_addr_out_reg[10] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_address [10]),
        .Q(\processor/wb_csr_address [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_addr_out_reg[11] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_address [11]),
        .Q(\processor/wb_csr_address [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_addr_out_reg[1] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_address [1]),
        .Q(\processor/wb_csr_address [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_addr_out_reg[2] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_address [2]),
        .Q(\processor/wb_csr_address [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_addr_out_reg[3] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_address [3]),
        .Q(\processor/wb_csr_address [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_addr_out_reg[4] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_address [4]),
        .Q(\processor/wb_csr_address [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_addr_out_reg[5] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_address [5]),
        .Q(\processor/wb_csr_address [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_addr_out_reg[6] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_address [6]),
        .Q(\processor/wb_csr_address [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_addr_out_reg[7] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_address [7]),
        .Q(\processor/wb_csr_address [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_addr_out_reg[8] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_address [8]),
        .Q(\processor/wb_csr_address [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_addr_out_reg[9] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_address [9]),
        .Q(\processor/wb_csr_address [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[0] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [0]),
        .Q(\processor/wb_csr_data [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[10] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [10]),
        .Q(\processor/wb_csr_data [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[11] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [11]),
        .Q(\processor/wb_csr_data [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[12] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [12]),
        .Q(\processor/wb_csr_data [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[13] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [13]),
        .Q(\processor/wb_csr_data [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[14] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [14]),
        .Q(\processor/wb_csr_data [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[15] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [15]),
        .Q(\processor/wb_csr_data [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[16] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [16]),
        .Q(\processor/wb_csr_data [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[17] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [17]),
        .Q(\processor/wb_csr_data [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[18] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [18]),
        .Q(\processor/wb_csr_data [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[19] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [19]),
        .Q(\processor/wb_csr_data [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[1] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [1]),
        .Q(\processor/wb_csr_data [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[20] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [20]),
        .Q(\processor/wb_csr_data [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[21] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [21]),
        .Q(\processor/wb_csr_data [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[22] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [22]),
        .Q(\processor/wb_csr_data [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[23] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [23]),
        .Q(\processor/wb_csr_data [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[24] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [24]),
        .Q(\processor/wb_csr_data [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[25] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [25]),
        .Q(\processor/wb_csr_data [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[26] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [26]),
        .Q(\processor/wb_csr_data [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[27] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [27]),
        .Q(\processor/wb_csr_data [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[28] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [28]),
        .Q(\processor/wb_csr_data [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[29] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [29]),
        .Q(\processor/wb_csr_data [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[2] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [2]),
        .Q(\processor/wb_csr_data [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[30] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [30]),
        .Q(\processor/wb_csr_data [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[31] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [31]),
        .Q(\processor/wb_csr_data [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[3] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [3]),
        .Q(\processor/wb_csr_data [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[4] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [4]),
        .Q(\processor/wb_csr_data [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[5] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [5]),
        .Q(\processor/wb_csr_data [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[6] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [6]),
        .Q(\processor/wb_csr_data [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[7] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [7]),
        .Q(\processor/wb_csr_data [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[8] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [8]),
        .Q(\processor/wb_csr_data [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_data_out_reg[9] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_data [9]),
        .Q(\processor/wb_csr_data [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_write_out_reg[0] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_write [0]),
        .Q(\processor/wb_csr_write [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/csr_write_out_reg[1] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_csr_write [1]),
        .Q(\processor/wb_csr_write [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][0] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [0]),
        .Q(\processor/wb_exception_context[badaddr] [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][10] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [10]),
        .Q(\processor/wb_exception_context[badaddr] [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][11] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [11]),
        .Q(\processor/wb_exception_context[badaddr] [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][12] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [12]),
        .Q(\processor/wb_exception_context[badaddr] [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][13] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [13]),
        .Q(\processor/wb_exception_context[badaddr] [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][14] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [14]),
        .Q(\processor/wb_exception_context[badaddr] [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][15] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [15]),
        .Q(\processor/wb_exception_context[badaddr] [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][16] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [16]),
        .Q(\processor/wb_exception_context[badaddr] [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][17] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [17]),
        .Q(\processor/wb_exception_context[badaddr] [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][18] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [18]),
        .Q(\processor/wb_exception_context[badaddr] [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][19] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [19]),
        .Q(\processor/wb_exception_context[badaddr] [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][1] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [1]),
        .Q(\processor/wb_exception_context[badaddr] [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][20] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [20]),
        .Q(\processor/wb_exception_context[badaddr] [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][21] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [21]),
        .Q(\processor/wb_exception_context[badaddr] [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][22] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [22]),
        .Q(\processor/wb_exception_context[badaddr] [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][23] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [23]),
        .Q(\processor/wb_exception_context[badaddr] [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][24] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [24]),
        .Q(\processor/wb_exception_context[badaddr] [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][25] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [25]),
        .Q(\processor/wb_exception_context[badaddr] [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][26] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [26]),
        .Q(\processor/wb_exception_context[badaddr] [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][27] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [27]),
        .Q(\processor/wb_exception_context[badaddr] [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][28] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [28]),
        .Q(\processor/wb_exception_context[badaddr] [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][29] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [29]),
        .Q(\processor/wb_exception_context[badaddr] [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][2] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [2]),
        .Q(\processor/wb_exception_context[badaddr] [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][30] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [30]),
        .Q(\processor/wb_exception_context[badaddr] [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][31] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [31]),
        .Q(\processor/wb_exception_context[badaddr] [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][3] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [3]),
        .Q(\processor/wb_exception_context[badaddr] [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][4] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [4]),
        .Q(\processor/wb_exception_context[badaddr] [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][5] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [5]),
        .Q(\processor/wb_exception_context[badaddr] [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][6] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [6]),
        .Q(\processor/wb_exception_context[badaddr] [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][7] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [7]),
        .Q(\processor/wb_exception_context[badaddr] [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][8] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [8]),
        .Q(\processor/wb_exception_context[badaddr] [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[badaddr][9] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[badaddr] [9]),
        .Q(\processor/wb_exception_context[badaddr] [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[cause][0] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[cause] [0]),
        .Q(\processor/wb_exception_context[cause] [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[cause][1] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[cause] [1]),
        .Q(\processor/wb_exception_context[cause] [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[cause][2] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[cause] [2]),
        .Q(\processor/wb_exception_context[cause] [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[cause][3] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[cause] [3]),
        .Q(\processor/wb_exception_context[cause] [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[cause][4] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[cause] [4]),
        .Q(\processor/wb_exception_context[cause] [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[cause][5] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[cause] [5]),
        .Q(\processor/wb_exception_context[cause] [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[ie1] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context ),
        .Q(\processor/wb_exception_context ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_ctx_out_reg[ie] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_exception_context[ie] ),
        .Q(\processor/wb_exception_context[ie] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/exception_out_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\processor/mem_exception ),
        .Q(\processor/wb_exception ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_addr_out_reg[0] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_address [0]),
        .Q(\processor/wb_rd_address [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_addr_out_reg[1] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_address [1]),
        .Q(\processor/wb_rd_address [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_addr_out_reg[2] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_address [2]),
        .Q(\processor/wb_rd_address [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_addr_out_reg[3] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_address [3]),
        .Q(\processor/wb_rd_address [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_addr_out_reg[4] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_address [4]),
        .Q(\processor/wb_rd_address [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[0] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_data [0]),
        .Q(\processor/wb_rd_data [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[10] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(rd_data_out),
        .Q(\processor/wb_rd_data [10]),
        .S(\rd_data_out[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[11] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\rd_data_out[11]_i_1_n_0 ),
        .Q(\processor/wb_rd_data [11]),
        .S(\rd_data_out[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[12] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\rd_data_out[12]_i_1_n_0 ),
        .Q(\processor/wb_rd_data [12]),
        .S(\rd_data_out[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[13] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\rd_data_out[13]_i_1_n_0 ),
        .Q(\processor/wb_rd_data [13]),
        .S(\rd_data_out[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[14] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\rd_data_out[14]_i_1_n_0 ),
        .Q(\processor/wb_rd_data [14]),
        .S(\rd_data_out[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[15] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\rd_data_out[15]_i_2_n_0 ),
        .Q(\processor/wb_rd_data [15]),
        .S(\rd_data_out[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[16] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_data [16]),
        .Q(\processor/wb_rd_data [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[17] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_data [17]),
        .Q(\processor/wb_rd_data [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[18] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_data [18]),
        .Q(\processor/wb_rd_data [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[19] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_data [19]),
        .Q(\processor/wb_rd_data [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[1] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_data [1]),
        .Q(\processor/wb_rd_data [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[20] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_data [20]),
        .Q(\processor/wb_rd_data [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[21] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_data [21]),
        .Q(\processor/wb_rd_data [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[22] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_data [22]),
        .Q(\processor/wb_rd_data [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[23] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_data [23]),
        .Q(\processor/wb_rd_data [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[24] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_data [24]),
        .Q(\processor/wb_rd_data [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[25] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_data [25]),
        .Q(\processor/wb_rd_data [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[26] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_data [26]),
        .Q(\processor/wb_rd_data [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[27] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_data [27]),
        .Q(\processor/wb_rd_data [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[28] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_data [28]),
        .Q(\processor/wb_rd_data [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[29] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_data [29]),
        .Q(\processor/wb_rd_data [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[2] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_data [2]),
        .Q(\processor/wb_rd_data [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[30] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_data [30]),
        .Q(\processor/wb_rd_data [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[31] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_data [31]),
        .Q(\processor/wb_rd_data [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[3] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_data [3]),
        .Q(\processor/wb_rd_data [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[4] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_data [4]),
        .Q(\processor/wb_rd_data [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[5] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_data [5]),
        .Q(\processor/wb_rd_data [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[6] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_data [6]),
        .Q(\processor/wb_rd_data [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[7] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\processor/mem_rd_data [7]),
        .Q(\processor/wb_rd_data [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[8] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\rd_data_out[8]_i_1_n_0 ),
        .Q(\processor/wb_rd_data [8]),
        .S(\rd_data_out[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \processor/writeback/rd_data_out_reg[9] 
       (.C(clk),
        .CE(\icache/p_3_in ),
        .D(\rd_data_out[9]_i_1_n_0 ),
        .Q(\processor/wb_rd_data [9]),
        .S(\rd_data_out[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \processor/writeback/rd_write_out_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\processor/mem_rd_write ),
        .Q(\processor/wb_rd_write ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rd_data[0]_i_11 
       (.I0(\rd_data[4]_i_11_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[0]_i_28_n_0 ),
        .I3(\processor/execute/alu_y [3]),
        .I4(\rd_data[0]_i_29_n_0 ),
        .O(\rd_data[0]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[0]_i_12 
       (.I0(\processor/execute/alu_x [24]),
        .I1(\processor/execute/alu_x [8]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_x [16]),
        .I4(\processor/execute/alu_y [4]),
        .I5(\processor/execute/alu_x [0]),
        .O(\rd_data[0]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \rd_data[0]_i_14 
       (.I0(\processor/execute/alu_y [30]),
        .I1(\processor/execute/alu_x [30]),
        .I2(\processor/execute/alu_x [31]),
        .I3(\processor/execute/alu_y [31]),
        .O(\rd_data[0]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \rd_data[0]_i_15 
       (.I0(\processor/execute/alu_y [28]),
        .I1(\processor/execute/alu_x [28]),
        .I2(\processor/execute/alu_x [29]),
        .I3(\processor/execute/alu_y [29]),
        .O(\rd_data[0]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \rd_data[0]_i_16 
       (.I0(\processor/execute/alu_y [26]),
        .I1(\processor/execute/alu_x [26]),
        .I2(\processor/execute/alu_x[27]_repN ),
        .I3(\processor/execute/alu_y [27]),
        .O(\rd_data[0]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \rd_data[0]_i_17 
       (.I0(\processor/execute/alu_y [24]),
        .I1(\processor/execute/alu_x [24]),
        .I2(\processor/execute/alu_x [25]),
        .I3(\processor/execute/alu_y [25]),
        .O(\rd_data[0]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_18 
       (.I0(\processor/execute/alu_x [30]),
        .I1(\processor/execute/alu_y [30]),
        .I2(\processor/execute/alu_x [31]),
        .I3(\processor/execute/alu_y [31]),
        .O(\rd_data[0]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_19 
       (.I0(\processor/execute/alu_x [28]),
        .I1(\processor/execute/alu_y [28]),
        .I2(\processor/execute/alu_x [29]),
        .I3(\processor/execute/alu_y [29]),
        .O(\rd_data[0]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[0]_i_2 
       (.I0(\rd_data[0]_i_4_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\rd_data[0]_i_5_n_0 ),
        .I3(\processor/execute/alu_op [2]),
        .I4(\rd_data[0]_i_6_n_0 ),
        .O(\rd_data[0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_20 
       (.I0(\processor/execute/alu_x [26]),
        .I1(\processor/execute/alu_y [26]),
        .I2(\processor/execute/alu_x[27]_repN ),
        .I3(\processor/execute/alu_y [27]),
        .O(\rd_data[0]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_21 
       (.I0(\processor/execute/alu_x [24]),
        .I1(\processor/execute/alu_y [24]),
        .I2(\processor/execute/alu_x [25]),
        .I3(\processor/execute/alu_y [25]),
        .O(\rd_data[0]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \rd_data[0]_i_23 
       (.I0(\processor/execute/alu_y [30]),
        .I1(\processor/execute/alu_x [30]),
        .I2(\processor/execute/alu_y [31]),
        .I3(\processor/execute/alu_x [31]),
        .O(\rd_data[0]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_24 
       (.I0(\processor/execute/alu_x [30]),
        .I1(\processor/execute/alu_y [30]),
        .I2(\processor/execute/alu_y [31]),
        .I3(\processor/execute/alu_x [31]),
        .O(\rd_data[0]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_25 
       (.I0(\processor/execute/alu_x [28]),
        .I1(\processor/execute/alu_y [28]),
        .I2(\processor/execute/alu_x [29]),
        .I3(\processor/execute/alu_y [29]),
        .O(\rd_data[0]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_26 
       (.I0(\processor/execute/alu_x [26]),
        .I1(\processor/execute/alu_y [26]),
        .I2(\processor/execute/alu_x[27]_repN ),
        .I3(\processor/execute/alu_y [27]),
        .O(\rd_data[0]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_27 
       (.I0(\processor/execute/alu_x [24]),
        .I1(\processor/execute/alu_y [24]),
        .I2(\processor/execute/alu_x [25]),
        .I3(\processor/execute/alu_y [25]),
        .O(\rd_data[0]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rd_data[0]_i_28 
       (.I0(\processor/execute/alu_x [24]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [8]),
        .O(\rd_data[0]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rd_data[0]_i_29 
       (.I0(\processor/execute/alu_x [16]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [0]),
        .O(\rd_data[0]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000F404)) 
    \rd_data[0]_i_3 
       (.I0(\processor/execute/alu_y [0]),
        .I1(\rd_data[1]_i_6_n_0 ),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data7 [0]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\processor/execute/alu_op [1]),
        .O(\rd_data[0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \rd_data[0]_i_31 
       (.I0(\processor/execute/alu_y [22]),
        .I1(\processor/execute/alu_x [22]),
        .I2(\processor/execute/alu_x [23]),
        .I3(\processor/execute/alu_y [23]),
        .O(\rd_data[0]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \rd_data[0]_i_32 
       (.I0(\processor/execute/alu_y [20]),
        .I1(\processor/execute/alu_x [20]),
        .I2(\processor/execute/alu_x [21]),
        .I3(\processor/execute/alu_y [21]),
        .O(\rd_data[0]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \rd_data[0]_i_33 
       (.I0(\processor/execute/alu_y [18]),
        .I1(\processor/execute/alu_x [18]),
        .I2(\processor/execute/alu_x [19]),
        .I3(\processor/execute/alu_y [19]),
        .O(\rd_data[0]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \rd_data[0]_i_34 
       (.I0(\processor/execute/alu_y [16]),
        .I1(\processor/execute/alu_x [16]),
        .I2(\processor/execute/alu_x [17]),
        .I3(\processor/execute/alu_y [17]),
        .O(\rd_data[0]_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_35 
       (.I0(\processor/execute/alu_x [22]),
        .I1(\processor/execute/alu_y [22]),
        .I2(\processor/execute/alu_x [23]),
        .I3(\processor/execute/alu_y [23]),
        .O(\rd_data[0]_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_36 
       (.I0(\processor/execute/alu_x [20]),
        .I1(\processor/execute/alu_y [20]),
        .I2(\processor/execute/alu_x [21]),
        .I3(\processor/execute/alu_y [21]),
        .O(\rd_data[0]_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_37 
       (.I0(\processor/execute/alu_x [18]),
        .I1(\processor/execute/alu_y [18]),
        .I2(\processor/execute/alu_x [19]),
        .I3(\processor/execute/alu_y [19]),
        .O(\rd_data[0]_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_38 
       (.I0(\processor/execute/alu_x [16]),
        .I1(\processor/execute/alu_y [16]),
        .I2(\processor/execute/alu_x [17]),
        .I3(\processor/execute/alu_y [17]),
        .O(\rd_data[0]_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[0]_i_4 
       (.I0(\rd_data[1]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[0]_i_8_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [0]),
        .O(\rd_data[0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_40 
       (.I0(\processor/execute/alu_x [22]),
        .I1(\processor/execute/alu_y [22]),
        .I2(\processor/execute/alu_x [23]),
        .I3(\processor/execute/alu_y [23]),
        .O(\rd_data[0]_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_41 
       (.I0(\processor/execute/alu_x [20]),
        .I1(\processor/execute/alu_y [20]),
        .I2(\processor/execute/alu_x [21]),
        .I3(\processor/execute/alu_y [21]),
        .O(\rd_data[0]_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_42 
       (.I0(\processor/execute/alu_x [18]),
        .I1(\processor/execute/alu_y [18]),
        .I2(\processor/execute/alu_x [19]),
        .I3(\processor/execute/alu_y [19]),
        .O(\rd_data[0]_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_43 
       (.I0(\processor/execute/alu_x [16]),
        .I1(\processor/execute/alu_y [16]),
        .I2(\processor/execute/alu_x [17]),
        .I3(\processor/execute/alu_y [17]),
        .O(\rd_data[0]_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \rd_data[0]_i_45 
       (.I0(\processor/execute/alu_y [14]),
        .I1(\processor/execute/alu_x [14]),
        .I2(\processor/execute/alu_x [15]),
        .I3(\processor/execute/alu_y [15]),
        .O(\rd_data[0]_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \rd_data[0]_i_46 
       (.I0(\processor/execute/alu_y [12]),
        .I1(\processor/execute/alu_x [12]),
        .I2(\processor/execute/alu_x [13]),
        .I3(\processor/execute/alu_y [13]),
        .O(\rd_data[0]_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \rd_data[0]_i_47 
       (.I0(\processor/execute/alu_y [10]),
        .I1(\processor/execute/alu_x [10]),
        .I2(\processor/execute/alu_x [11]),
        .I3(\processor/execute/alu_y [11]),
        .O(\rd_data[0]_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \rd_data[0]_i_48 
       (.I0(\processor/execute/alu_y [8]),
        .I1(\processor/execute/alu_x [8]),
        .I2(\processor/execute/alu_x [9]),
        .I3(\processor/execute/alu_y [9]),
        .O(\rd_data[0]_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_49 
       (.I0(\processor/execute/alu_x [14]),
        .I1(\processor/execute/alu_y [14]),
        .I2(\processor/execute/alu_x [15]),
        .I3(\processor/execute/alu_y [15]),
        .O(\rd_data[0]_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rd_data[0]_i_5 
       (.I0(\processor/execute/alu_instance/data5 [0]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_instance/data4 ),
        .O(\rd_data[0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_50 
       (.I0(\processor/execute/alu_x [12]),
        .I1(\processor/execute/alu_y [12]),
        .I2(\processor/execute/alu_x [13]),
        .I3(\processor/execute/alu_y [13]),
        .O(\rd_data[0]_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_51 
       (.I0(\processor/execute/alu_x [10]),
        .I1(\processor/execute/alu_y [10]),
        .I2(\processor/execute/alu_x [11]),
        .I3(\processor/execute/alu_y [11]),
        .O(\rd_data[0]_i_51_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_52 
       (.I0(\processor/execute/alu_x [8]),
        .I1(\processor/execute/alu_y [8]),
        .I2(\processor/execute/alu_x [9]),
        .I3(\processor/execute/alu_y [9]),
        .O(\rd_data[0]_i_52_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_54 
       (.I0(\processor/execute/alu_x [14]),
        .I1(\processor/execute/alu_y [14]),
        .I2(\processor/execute/alu_x [15]),
        .I3(\processor/execute/alu_y [15]),
        .O(\rd_data[0]_i_54_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_55 
       (.I0(\processor/execute/alu_x [12]),
        .I1(\processor/execute/alu_y [12]),
        .I2(\processor/execute/alu_x [13]),
        .I3(\processor/execute/alu_y [13]),
        .O(\rd_data[0]_i_55_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_56 
       (.I0(\processor/execute/alu_x [10]),
        .I1(\processor/execute/alu_y [10]),
        .I2(\processor/execute/alu_x [11]),
        .I3(\processor/execute/alu_y [11]),
        .O(\rd_data[0]_i_56_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_57 
       (.I0(\processor/execute/alu_x [8]),
        .I1(\processor/execute/alu_y [8]),
        .I2(\processor/execute/alu_x [9]),
        .I3(\processor/execute/alu_y [9]),
        .O(\rd_data[0]_i_57_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \rd_data[0]_i_58 
       (.I0(\processor/execute/alu_y [6]),
        .I1(\processor/execute/alu_x [6]),
        .I2(\processor/execute/alu_x [7]),
        .I3(\processor/execute/alu_y [7]),
        .O(\rd_data[0]_i_58_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \rd_data[0]_i_59 
       (.I0(\processor/execute/alu_y [4]),
        .I1(\processor/execute/alu_x [4]),
        .I2(\processor/execute/alu_x [5]),
        .I3(\processor/execute/alu_y [5]),
        .O(\rd_data[0]_i_59_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB3BCBC80)) 
    \rd_data[0]_i_6 
       (.I0(\processor/execute/alu_instance/data3 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_x [0]),
        .I4(\processor/execute/alu_y [0]),
        .O(\rd_data[0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \rd_data[0]_i_60 
       (.I0(\processor/execute/alu_y [2]),
        .I1(\processor/execute/alu_x [2]),
        .I2(\processor/execute/alu_x [3]),
        .I3(\processor/execute/alu_y [3]),
        .O(\rd_data[0]_i_60_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \rd_data[0]_i_61 
       (.I0(\processor/execute/alu_y [0]),
        .I1(\processor/execute/alu_x [0]),
        .I2(\processor/execute/alu_x [1]),
        .I3(\processor/execute/alu_y [1]),
        .O(\rd_data[0]_i_61_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_62 
       (.I0(\processor/execute/alu_x [6]),
        .I1(\processor/execute/alu_y [6]),
        .I2(\processor/execute/alu_x [7]),
        .I3(\processor/execute/alu_y [7]),
        .O(\rd_data[0]_i_62_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_63 
       (.I0(\processor/execute/alu_x [4]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [5]),
        .I3(\processor/execute/alu_y [5]),
        .O(\rd_data[0]_i_63_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_64 
       (.I0(\processor/execute/alu_x [2]),
        .I1(\processor/execute/alu_y [2]),
        .I2(\processor/execute/alu_x [3]),
        .I3(\processor/execute/alu_y [3]),
        .O(\rd_data[0]_i_64_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_65 
       (.I0(\processor/execute/alu_x [1]),
        .I1(\processor/execute/alu_y [1]),
        .I2(\processor/execute/alu_x [0]),
        .I3(\processor/execute/alu_y [0]),
        .O(\rd_data[0]_i_65_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_66 
       (.I0(\processor/execute/alu_x [6]),
        .I1(\processor/execute/alu_y [6]),
        .I2(\processor/execute/alu_x [7]),
        .I3(\processor/execute/alu_y [7]),
        .O(\rd_data[0]_i_66_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_67 
       (.I0(\processor/execute/alu_x [4]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [5]),
        .I3(\processor/execute/alu_y [5]),
        .O(\rd_data[0]_i_67_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_68 
       (.I0(\processor/execute/alu_x [2]),
        .I1(\processor/execute/alu_y [2]),
        .I2(\processor/execute/alu_x [3]),
        .I3(\processor/execute/alu_y [3]),
        .O(\rd_data[0]_i_68_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \rd_data[0]_i_69 
       (.I0(\processor/execute/alu_x [1]),
        .I1(\processor/execute/alu_y [1]),
        .I2(\processor/execute/alu_x [0]),
        .I3(\processor/execute/alu_y [0]),
        .O(\rd_data[0]_i_69_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rd_data[0]_i_7 
       (.I0(\rd_data[1]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[2]_i_14_n_0 ),
        .I3(\processor/execute/alu_y [1]),
        .I4(\rd_data[0]_i_11_n_0 ),
        .O(\processor/execute/alu_instance/data7 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[0]_i_8 
       (.I0(\rd_data[6]_i_8_n_0 ),
        .I1(\rd_data[1]_i_10_n_0 ),
        .I2(\processor/execute/alu_y [1]),
        .I3(\rd_data[4]_i_11_n_0 ),
        .I4(\processor/execute/alu_y [2]),
        .I5(\rd_data[0]_i_12_n_0 ),
        .O(\rd_data[0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[10]_i_1 
       (.I0(\rd_data[10]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[10]_i_3_n_0 ),
        .O(\processor/ex_rd_data [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[10]_i_10 
       (.I0(\rd_data[16]_i_13_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[12]_i_12_n_0 ),
        .I3(\rd_data[14]_i_12_n_0 ),
        .I4(\rd_data[10]_i_13_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[10]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[10]_i_11 
       (.I0(\rd_data[10]_i_14_n_0 ),
        .I1(\csr_data_out[10]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [10]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rd_data[10]_i_12 
       (.I0(\processor/execute/alu_x [26]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [10]),
        .O(\rd_data[10]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \rd_data[10]_i_13 
       (.I0(\processor/execute/alu_x [18]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\rd_data[10]_i_12_n_0 ),
        .O(\rd_data[10]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[10]_i_14 
       (.I0(\processor/ex_pc [10]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [10]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [10]),
        .O(\rd_data[10]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[10]_i_2 
       (.I0(\rd_data[11]_i_4_n_0 ),
        .I1(\rd_data[10]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[10]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[11]_i_5_n_0 ),
        .O(\rd_data[10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[10]_i_3 
       (.I0(\rd_data[10]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [10]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[10]_i_7_n_0 ),
        .O(\rd_data[10]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[10]_i_4 
       (.I0(\rd_data[14]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[10]_i_8_n_0 ),
        .I3(\rd_data[16]_i_8_n_0 ),
        .I4(\rd_data[12]_i_8_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[10]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[10]_i_5 
       (.I0(\rd_data[10]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[14]_i_9_n_0 ),
        .I3(\rd_data[12]_i_9_n_0 ),
        .I4(\rd_data[16]_i_9_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[10]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[10]_i_6 
       (.I0(\rd_data[11]_i_11_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[10]_i_10_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [10]),
        .O(\rd_data[10]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[10]_i_7 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [10]),
        .I3(\processor/execute/alu_y [10]),
        .O(\rd_data[10]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[10]_i_8 
       (.I0(\processor/execute/alu_x [31]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [18]),
        .I3(\processor/execute/alu_y [3]),
        .I4(\rd_data[10]_i_12_n_0 ),
        .O(\rd_data[10]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \rd_data[10]_i_9 
       (.I0(\processor/execute/alu_x [3]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_y [3]),
        .O(\rd_data[10]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[11]_i_1 
       (.I0(\rd_data[11]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[11]_i_3_n_0 ),
        .O(\processor/ex_rd_data [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h04FF0400)) 
    \rd_data[11]_i_10 
       (.I0(\processor/execute/alu_y [4]),
        .I1(\processor/execute/alu_x [4]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_y [2]),
        .I4(\rd_data[15]_i_10_n_0 ),
        .O(\rd_data[11]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[11]_i_11 
       (.I0(\rd_data[17]_i_13_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[13]_i_12_n_0 ),
        .I3(\rd_data[15]_i_22_n_0 ),
        .I4(\rd_data[11]_i_23_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[11]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[11]_i_13 
       (.I0(\rd_data[11]_i_28_n_0 ),
        .I1(\rd_data[11]_i_29_n_0 ),
        .I2(\rd_data[11]_i_30_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [11]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[11]_i_14 
       (.I0(\rd_data[11]_i_31_n_0 ),
        .I1(\rd_data[11]_i_32_n_0 ),
        .I2(\rd_data[11]_i_33_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [10]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[11]_i_15 
       (.I0(\rd_data[11]_i_34_n_0 ),
        .I1(\rd_data[11]_i_35_n_0 ),
        .I2(\rd_data[11]_i_36_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [9]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[11]_i_16 
       (.I0(\rd_data[11]_i_37_n_0 ),
        .I1(\rd_data[11]_i_38_n_0 ),
        .I2(\rd_data[11]_i_39_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [8]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[11]_i_17 
       (.I0(\processor/execute/alu_x [11]),
        .I1(\processor/execute/alu_y [11]),
        .O(\rd_data[11]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[11]_i_18 
       (.I0(\processor/execute/alu_x [10]),
        .I1(\processor/execute/alu_y [10]),
        .O(\rd_data[11]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[11]_i_19 
       (.I0(\processor/execute/alu_x [9]),
        .I1(\processor/execute/alu_y [9]),
        .O(\rd_data[11]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[11]_i_2 
       (.I0(\rd_data[12]_i_4_n_0 ),
        .I1(\rd_data[11]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[11]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[12]_i_5_n_0 ),
        .O(\rd_data[11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[11]_i_20 
       (.I0(\processor/execute/alu_x [8]),
        .I1(\processor/execute/alu_y [8]),
        .O(\rd_data[11]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[11]_i_21 
       (.I0(\rd_data[11]_i_41_n_0 ),
        .I1(\csr_data_out[11]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [11]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rd_data[11]_i_22 
       (.I0(\processor/execute/alu_x [27]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [11]),
        .O(\rd_data[11]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \rd_data[11]_i_23 
       (.I0(\processor/execute/alu_x [19]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\rd_data[11]_i_22_n_0 ),
        .O(\rd_data[11]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[11]_i_24 
       (.I0(\processor/execute/alu_x [11]),
        .I1(\processor/execute/alu_y [11]),
        .O(\rd_data[11]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[11]_i_25 
       (.I0(\processor/execute/alu_x [10]),
        .I1(\processor/execute/alu_y [10]),
        .O(\rd_data[11]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[11]_i_26 
       (.I0(\processor/execute/alu_x [9]),
        .I1(\processor/execute/alu_y [9]),
        .O(\rd_data[11]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[11]_i_27 
       (.I0(\processor/execute/alu_x [8]),
        .I1(\processor/execute/alu_y [8]),
        .O(\rd_data[11]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[11]_i_28 
       (.I0(\processor/ex_pc [11]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [11]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [11]),
        .O(\rd_data[11]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \rd_data[11]_i_29 
       (.I0(\csr_data_out[11]_i_7_n_0 ),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [11]),
        .O(\rd_data[11]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[11]_i_3 
       (.I0(\rd_data[11]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [11]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[11]_i_8_n_0 ),
        .O(\rd_data[11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4545454444444544)) 
    \rd_data[11]_i_30 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\csr_data_out[11]_i_6_n_0 ),
        .I2(\csr_data_out[4]_i_9_n_0 ),
        .I3(\rd_data[11]_i_42_n_0 ),
        .I4(\csr_data_out[30]_i_9_n_0 ),
        .I5(\processor/wb_exception_context[badaddr] [11]),
        .O(\rd_data[11]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[11]_i_31 
       (.I0(\processor/ex_pc [10]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [10]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [10]),
        .O(\rd_data[11]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \rd_data[11]_i_32 
       (.I0(\csr_data_out[11]_i_7_n_0 ),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [10]),
        .O(\rd_data[11]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4545454444444544)) 
    \rd_data[11]_i_33 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\csr_data_out[10]_i_6_n_0 ),
        .I2(\csr_data_out[4]_i_9_n_0 ),
        .I3(\rd_data[11]_i_43_n_0 ),
        .I4(\csr_data_out[30]_i_9_n_0 ),
        .I5(\processor/wb_exception_context[badaddr] [10]),
        .O(\rd_data[11]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[11]_i_34 
       (.I0(\processor/ex_pc [9]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [9]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [9]),
        .O(\rd_data[11]_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rd_data[11]_i_35 
       (.I0(\processor/mem_exception_context[badaddr] [9]),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .O(\rd_data[11]_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000540455555555)) 
    \rd_data[11]_i_36 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\rd_data[11]_i_44_n_0 ),
        .I2(\csr_data_out[30]_i_9_n_0 ),
        .I3(\processor/wb_exception_context[badaddr] [9]),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\rd_data[11]_i_45_n_0 ),
        .O(\rd_data[11]_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[11]_i_37 
       (.I0(\processor/ex_pc [8]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [8]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [8]),
        .O(\rd_data[11]_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \rd_data[11]_i_38 
       (.I0(\csr_data_out[11]_i_7_n_0 ),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [8]),
        .O(\rd_data[11]_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4545454444444544)) 
    \rd_data[11]_i_39 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\csr_data_out[8]_i_6_n_0 ),
        .I2(\csr_data_out[4]_i_9_n_0 ),
        .I3(\rd_data[11]_i_46_n_0 ),
        .I4(\csr_data_out[30]_i_9_n_0 ),
        .I5(\processor/wb_exception_context[badaddr] [8]),
        .O(\rd_data[11]_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[11]_i_4 
       (.I0(\rd_data[17]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[13]_i_8_n_0 ),
        .I3(\rd_data[15]_i_9_n_0 ),
        .I4(\rd_data[11]_i_9_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[11]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[11]_i_41 
       (.I0(\processor/ex_pc [11]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [11]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [11]),
        .O(\rd_data[11]_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEAEAEAAA2A2A2AAA)) 
    \rd_data[11]_i_42 
       (.I0(\processor/csr_read_data [11]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded3 ),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/wb_csr_write [0]),
        .I5(\processor/wb_csr_data [11]),
        .O(\rd_data[11]_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEAEAEAAA2A2A2AAA)) 
    \rd_data[11]_i_43 
       (.I0(\processor/csr_read_data [10]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded3 ),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/wb_csr_write [0]),
        .I5(\processor/wb_csr_data [10]),
        .O(\rd_data[11]_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCAAACAAACAAAAAAA)) 
    \rd_data[11]_i_44 
       (.I0(\processor/csr_read_data [9]),
        .I1(\processor/wb_csr_data [9]),
        .I2(\processor/execute/csr_writeable ),
        .I3(\processor/execute/csr_value_forwarded3 ),
        .I4(\processor/wb_csr_write [1]),
        .I5(\processor/wb_csr_write [0]),
        .O(\rd_data[11]_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7F7F7FFF)) 
    \rd_data[11]_i_45 
       (.I0(\processor/mem_csr_data [9]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/mem_csr_write [0]),
        .I4(\processor/mem_csr_write [1]),
        .O(\rd_data[11]_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEAEAEAAA2A2A2AAA)) 
    \rd_data[11]_i_46 
       (.I0(\processor/csr_read_data [8]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded3 ),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/wb_csr_write [0]),
        .I5(\processor/wb_csr_data [8]),
        .O(\rd_data[11]_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \rd_data[11]_i_5 
       (.I0(\rd_data[13]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[17]_i_9_n_0 ),
        .I3(\rd_data[11]_i_10_n_0 ),
        .I4(\processor/execute/alu_y [1]),
        .O(\rd_data[11]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[11]_i_6 
       (.I0(\rd_data[12]_i_10_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[11]_i_11_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [11]),
        .O(\rd_data[11]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[11]_i_8 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [11]),
        .I3(\processor/execute/alu_y [11]),
        .O(\rd_data[11]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[11]_i_9 
       (.I0(\processor/execute/alu_x [31]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [19]),
        .I3(\processor/execute/alu_y [3]),
        .I4(\rd_data[11]_i_22_n_0 ),
        .O(\rd_data[11]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[12]_i_1 
       (.I0(\rd_data[12]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[12]_i_3_n_0 ),
        .O(\processor/ex_rd_data [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[12]_i_10 
       (.I0(\rd_data[16]_i_13_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[12]_i_12_n_0 ),
        .I3(\rd_data[18]_i_13_n_0 ),
        .I4(\rd_data[14]_i_12_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[12]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[12]_i_11 
       (.I0(\rd_data[12]_i_13_n_0 ),
        .I1(\csr_data_out[12]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [12]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h3300B8B8)) 
    \rd_data[12]_i_12 
       (.I0(\processor/execute/alu_x [28]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [12]),
        .I3(\processor/execute/alu_x [20]),
        .I4(\processor/execute/alu_y [3]),
        .O(\rd_data[12]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[12]_i_13 
       (.I0(\processor/ex_pc [12]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [12]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [12]),
        .O(\rd_data[12]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[12]_i_2 
       (.I0(\rd_data[13]_i_4_n_0 ),
        .I1(\rd_data[12]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[12]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[13]_i_5_n_0 ),
        .O(\rd_data[12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[12]_i_3 
       (.I0(\rd_data[12]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [12]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[12]_i_7_n_0 ),
        .O(\rd_data[12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[12]_i_4 
       (.I0(\rd_data[16]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[12]_i_8_n_0 ),
        .I3(\rd_data[18]_i_8_n_0 ),
        .I4(\rd_data[14]_i_8_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[12]_i_5 
       (.I0(\rd_data[12]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[16]_i_9_n_0 ),
        .I3(\rd_data[14]_i_9_n_0 ),
        .I4(\rd_data[18]_i_9_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[12]_i_6 
       (.I0(\rd_data[13]_i_10_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[12]_i_10_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [12]),
        .O(\rd_data[12]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[12]_i_7 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [12]),
        .I3(\processor/execute/alu_y [12]),
        .O(\rd_data[12]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[12]_i_8 
       (.I0(\processor/execute/alu_x [28]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [12]),
        .I3(\processor/execute/alu_x [31]),
        .I4(\processor/execute/alu_x [20]),
        .I5(\processor/execute/alu_y [3]),
        .O(\rd_data[12]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \rd_data[12]_i_9 
       (.I0(\processor/execute/alu_y [4]),
        .I1(\processor/execute/alu_x [5]),
        .I2(\processor/execute/alu_y [3]),
        .O(\rd_data[12]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[13]_i_1 
       (.I0(\rd_data[13]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[13]_i_3_n_0 ),
        .O(\processor/ex_rd_data [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[13]_i_10 
       (.I0(\rd_data[17]_i_13_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[13]_i_12_n_0 ),
        .I3(\rd_data[19]_i_24_n_0 ),
        .I4(\rd_data[15]_i_22_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[13]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[13]_i_11 
       (.I0(\rd_data[13]_i_13_n_0 ),
        .I1(\csr_data_out[13]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [13]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h3300B8B8)) 
    \rd_data[13]_i_12 
       (.I0(\processor/execute/alu_x [29]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [13]),
        .I3(\processor/execute/alu_x [21]),
        .I4(\processor/execute/alu_y [3]),
        .O(\rd_data[13]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[13]_i_13 
       (.I0(\processor/ex_pc [13]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [13]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [13]),
        .O(\rd_data[13]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[13]_i_2 
       (.I0(\rd_data[14]_i_4_n_0 ),
        .I1(\rd_data[13]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[13]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[14]_i_5_n_0 ),
        .O(\rd_data[13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[13]_i_3 
       (.I0(\rd_data[13]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [13]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[13]_i_7_n_0 ),
        .O(\rd_data[13]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[13]_i_4 
       (.I0(\rd_data[17]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[13]_i_8_n_0 ),
        .I3(\rd_data[19]_i_10_n_0 ),
        .I4(\rd_data[15]_i_9_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[13]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[13]_i_5 
       (.I0(\rd_data[13]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[17]_i_9_n_0 ),
        .I3(\rd_data[15]_i_10_n_0 ),
        .I4(\rd_data[19]_i_11_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[13]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[13]_i_6 
       (.I0(\rd_data[14]_i_10_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[13]_i_10_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [13]),
        .O(\rd_data[13]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[13]_i_7 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [13]),
        .I3(\processor/execute/alu_y [13]),
        .O(\rd_data[13]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[13]_i_8 
       (.I0(\processor/execute/alu_x [29]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [13]),
        .I3(\processor/execute/alu_x [31]),
        .I4(\processor/execute/alu_x [21]),
        .I5(\processor/execute/alu_y [3]),
        .O(\rd_data[13]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \rd_data[13]_i_9 
       (.I0(\processor/execute/alu_y [4]),
        .I1(\processor/execute/alu_x [6]),
        .I2(\processor/execute/alu_y [3]),
        .O(\rd_data[13]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[14]_i_1 
       (.I0(\rd_data[14]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[14]_i_3_n_0 ),
        .O(\processor/ex_rd_data [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[14]_i_10 
       (.I0(\rd_data[16]_i_12_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[16]_i_13_n_0 ),
        .I3(\rd_data[18]_i_13_n_0 ),
        .I4(\rd_data[14]_i_12_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[14]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[14]_i_11 
       (.I0(\rd_data[14]_i_13_n_0 ),
        .I1(\csr_data_out[14]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [14]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h3300B8B8)) 
    \rd_data[14]_i_12 
       (.I0(\processor/execute/alu_x [30]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [14]),
        .I3(\processor/execute/alu_x [22]),
        .I4(\processor/execute/alu_y [3]),
        .O(\rd_data[14]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[14]_i_13 
       (.I0(\processor/ex_pc [14]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [14]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [14]),
        .O(\rd_data[14]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[14]_i_2 
       (.I0(\rd_data[15]_i_4_n_0 ),
        .I1(\rd_data[14]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[14]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[15]_i_5_n_0 ),
        .O(\rd_data[14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[14]_i_3 
       (.I0(\rd_data[14]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [14]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[14]_i_7_n_0 ),
        .O(\rd_data[14]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[14]_i_4 
       (.I0(\rd_data[18]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[14]_i_8_n_0 ),
        .I3(\rd_data[20]_i_9_n_0 ),
        .I4(\rd_data[16]_i_8_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[14]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[14]_i_5 
       (.I0(\rd_data[14]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[18]_i_9_n_0 ),
        .I3(\rd_data[16]_i_9_n_0 ),
        .I4(\rd_data[20]_i_10_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[14]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[14]_i_6 
       (.I0(\rd_data[15]_i_11_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[14]_i_10_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [14]),
        .O(\rd_data[14]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[14]_i_7 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [14]),
        .I3(\processor/execute/alu_y [14]),
        .O(\rd_data[14]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[14]_i_8 
       (.I0(\processor/execute/alu_x [30]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [14]),
        .I3(\processor/execute/alu_x [31]),
        .I4(\processor/execute/alu_x [22]),
        .I5(\processor/execute/alu_y [3]),
        .O(\rd_data[14]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \rd_data[14]_i_9 
       (.I0(\processor/execute/alu_y [4]),
        .I1(\processor/execute/alu_x [7]),
        .I2(\processor/execute/alu_y [3]),
        .O(\rd_data[14]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[15]_i_1 
       (.I0(\rd_data[15]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[15]_i_3_n_0 ),
        .O(\processor/ex_rd_data [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2320)) 
    \rd_data[15]_i_10 
       (.I0(\processor/execute/alu_x [0]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_x [8]),
        .O(\rd_data[15]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[15]_i_11 
       (.I0(\rd_data[17]_i_12_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[17]_i_13_n_0 ),
        .I3(\rd_data[19]_i_24_n_0 ),
        .I4(\rd_data[15]_i_22_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[15]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[15]_i_13 
       (.I0(\rd_data[15]_i_27_n_0 ),
        .I1(\rd_data[15]_i_28_n_0 ),
        .I2(\rd_data[15]_i_29_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [15]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[15]_i_14 
       (.I0(\rd_data[15]_i_30_n_0 ),
        .I1(\rd_data[15]_i_31_n_0 ),
        .I2(\rd_data[15]_i_32_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [14]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[15]_i_15 
       (.I0(\rd_data[15]_i_33_n_0 ),
        .I1(\rd_data[15]_i_34_n_0 ),
        .I2(\rd_data[15]_i_35_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [13]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[15]_i_16 
       (.I0(\rd_data[15]_i_36_n_0 ),
        .I1(\rd_data[15]_i_37_n_0 ),
        .I2(\rd_data[15]_i_38_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [12]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[15]_i_17 
       (.I0(\processor/execute/alu_x [15]),
        .I1(\processor/execute/alu_y [15]),
        .O(\rd_data[15]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[15]_i_18 
       (.I0(\processor/execute/alu_x [14]),
        .I1(\processor/execute/alu_y [14]),
        .O(\rd_data[15]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[15]_i_19 
       (.I0(\processor/execute/alu_x [13]),
        .I1(\processor/execute/alu_y [13]),
        .O(\rd_data[15]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[15]_i_2 
       (.I0(\rd_data[16]_i_4_n_0 ),
        .I1(\rd_data[15]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[15]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[16]_i_5_n_0 ),
        .O(\rd_data[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[15]_i_20 
       (.I0(\processor/execute/alu_x [12]),
        .I1(\processor/execute/alu_y [12]),
        .O(\rd_data[15]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[15]_i_21 
       (.I0(\rd_data[15]_i_40_n_0 ),
        .I1(\csr_data_out[15]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [15]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h3300B8B8)) 
    \rd_data[15]_i_22 
       (.I0(\processor/execute/alu_x [31]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [15]),
        .I3(\processor/execute/alu_x [23]),
        .I4(\processor/execute/alu_y [3]),
        .O(\rd_data[15]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[15]_i_23 
       (.I0(\processor/execute/alu_x [15]),
        .I1(\processor/execute/alu_y [15]),
        .O(\rd_data[15]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[15]_i_24 
       (.I0(\processor/execute/alu_x [14]),
        .I1(\processor/execute/alu_y [14]),
        .O(\rd_data[15]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[15]_i_25 
       (.I0(\processor/execute/alu_x [13]),
        .I1(\processor/execute/alu_y [13]),
        .O(\rd_data[15]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[15]_i_26 
       (.I0(\processor/execute/alu_x [12]),
        .I1(\processor/execute/alu_y [12]),
        .O(\rd_data[15]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[15]_i_27 
       (.I0(\processor/ex_pc [15]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [15]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [15]),
        .O(\rd_data[15]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rd_data[15]_i_28 
       (.I0(\processor/mem_exception_context[badaddr] [15]),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .O(\rd_data[15]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000540455555555)) 
    \rd_data[15]_i_29 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\rd_data[15]_i_41_n_0 ),
        .I2(\csr_data_out[30]_i_9_n_0 ),
        .I3(\processor/wb_exception_context[badaddr] [15]),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\rd_data[15]_i_42_n_0 ),
        .O(\rd_data[15]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[15]_i_3 
       (.I0(\rd_data[15]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [15]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[15]_i_8_n_0 ),
        .O(\rd_data[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[15]_i_30 
       (.I0(\processor/ex_pc [14]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [14]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [14]),
        .O(\rd_data[15]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rd_data[15]_i_31 
       (.I0(\processor/mem_exception_context[badaddr] [14]),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .O(\rd_data[15]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000540455555555)) 
    \rd_data[15]_i_32 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\rd_data[15]_i_43_n_0 ),
        .I2(\csr_data_out[30]_i_9_n_0 ),
        .I3(\processor/wb_exception_context[badaddr] [14]),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\rd_data[15]_i_44_n_0 ),
        .O(\rd_data[15]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[15]_i_33 
       (.I0(\processor/ex_pc [13]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [13]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [13]),
        .O(\rd_data[15]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rd_data[15]_i_34 
       (.I0(\processor/mem_exception_context[badaddr] [13]),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .O(\rd_data[15]_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000540455555555)) 
    \rd_data[15]_i_35 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\rd_data[15]_i_45_n_0 ),
        .I2(\csr_data_out[30]_i_9_n_0 ),
        .I3(\processor/wb_exception_context[badaddr] [13]),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\rd_data[15]_i_46_n_0 ),
        .O(\rd_data[15]_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[15]_i_36 
       (.I0(\processor/ex_pc [12]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [12]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [12]),
        .O(\rd_data[15]_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rd_data[15]_i_37 
       (.I0(\processor/mem_exception_context[badaddr] [12]),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .O(\rd_data[15]_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000540455555555)) 
    \rd_data[15]_i_38 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\rd_data[15]_i_47_n_0 ),
        .I2(\csr_data_out[30]_i_9_n_0 ),
        .I3(\processor/wb_exception_context[badaddr] [12]),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\rd_data[15]_i_48_n_0 ),
        .O(\rd_data[15]_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[15]_i_4 
       (.I0(\rd_data[21]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[17]_i_8_n_0 ),
        .I3(\rd_data[19]_i_10_n_0 ),
        .I4(\rd_data[15]_i_9_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[15]_i_40 
       (.I0(\processor/ex_pc [15]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [15]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [15]),
        .O(\rd_data[15]_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCAAACAAACAAAAAAA)) 
    \rd_data[15]_i_41 
       (.I0(\processor/csr_read_data [15]),
        .I1(\processor/wb_csr_data [15]),
        .I2(\processor/execute/csr_writeable ),
        .I3(\processor/execute/csr_value_forwarded3 ),
        .I4(\processor/wb_csr_write [1]),
        .I5(\processor/wb_csr_write [0]),
        .O(\rd_data[15]_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7F7F7FFF)) 
    \rd_data[15]_i_42 
       (.I0(\processor/mem_csr_data [15]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/mem_csr_write [0]),
        .I4(\processor/mem_csr_write [1]),
        .O(\rd_data[15]_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCAAACAAACAAAAAAA)) 
    \rd_data[15]_i_43 
       (.I0(\processor/csr_read_data [14]),
        .I1(\processor/wb_csr_data [14]),
        .I2(\processor/execute/csr_writeable ),
        .I3(\processor/execute/csr_value_forwarded3 ),
        .I4(\processor/wb_csr_write [1]),
        .I5(\processor/wb_csr_write [0]),
        .O(\rd_data[15]_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7F7F7FFF)) 
    \rd_data[15]_i_44 
       (.I0(\processor/mem_csr_data [14]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/mem_csr_write [0]),
        .I4(\processor/mem_csr_write [1]),
        .O(\rd_data[15]_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCAAACAAACAAAAAAA)) 
    \rd_data[15]_i_45 
       (.I0(\processor/csr_read_data [13]),
        .I1(\processor/wb_csr_data [13]),
        .I2(\processor/execute/csr_writeable ),
        .I3(\processor/execute/csr_value_forwarded3 ),
        .I4(\processor/wb_csr_write [1]),
        .I5(\processor/wb_csr_write [0]),
        .O(\rd_data[15]_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7F7F7FFF)) 
    \rd_data[15]_i_46 
       (.I0(\processor/mem_csr_data [13]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/mem_csr_write [0]),
        .I4(\processor/mem_csr_write [1]),
        .O(\rd_data[15]_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCAAACAAACAAAAAAA)) 
    \rd_data[15]_i_47 
       (.I0(\processor/csr_read_data [12]),
        .I1(\processor/wb_csr_data [12]),
        .I2(\processor/execute/csr_writeable ),
        .I3(\processor/execute/csr_value_forwarded3 ),
        .I4(\processor/wb_csr_write [1]),
        .I5(\processor/wb_csr_write [0]),
        .O(\rd_data[15]_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7F7F7FFF)) 
    \rd_data[15]_i_48 
       (.I0(\processor/mem_csr_data [12]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/mem_csr_write [0]),
        .I4(\processor/mem_csr_write [1]),
        .O(\rd_data[15]_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[15]_i_5 
       (.I0(\rd_data[17]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[21]_i_10_n_0 ),
        .I3(\rd_data[15]_i_10_n_0 ),
        .I4(\rd_data[19]_i_11_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[15]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[15]_i_6 
       (.I0(\rd_data[16]_i_10_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[15]_i_11_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [15]),
        .O(\rd_data[15]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[15]_i_8 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [15]),
        .I3(\processor/execute/alu_y [15]),
        .O(\rd_data[15]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBB88B8B8)) 
    \rd_data[15]_i_9 
       (.I0(\processor/execute/alu_x [31]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [15]),
        .I3(\processor/execute/alu_x [23]),
        .I4(\processor/execute/alu_y [3]),
        .O(\rd_data[15]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[16]_i_1 
       (.I0(\rd_data[16]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[16]_i_3_n_0 ),
        .O(\processor/ex_rd_data [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[16]_i_10 
       (.I0(\rd_data[16]_i_12_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[16]_i_13_n_0 ),
        .I3(\rd_data[18]_i_12_n_0 ),
        .I4(\rd_data[18]_i_13_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[16]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[16]_i_11 
       (.I0(\rd_data[16]_i_14_n_0 ),
        .I1(\csr_data_out[16]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [16]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \rd_data[16]_i_12 
       (.I0(\processor/execute/alu_x [28]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [20]),
        .I3(\processor/execute/alu_y [4]),
        .O(\rd_data[16]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \rd_data[16]_i_13 
       (.I0(\processor/execute/alu_x [24]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [16]),
        .I3(\processor/execute/alu_y [4]),
        .O(\rd_data[16]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[16]_i_14 
       (.I0(\processor/ex_pc [16]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [16]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [16]),
        .O(\rd_data[16]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[16]_i_2 
       (.I0(\rd_data[17]_i_4_n_0 ),
        .I1(\rd_data[16]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[16]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[17]_i_5_n_0 ),
        .O(\rd_data[16]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[16]_i_3 
       (.I0(\rd_data[16]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [16]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[16]_i_7_n_0 ),
        .O(\rd_data[16]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[16]_i_4 
       (.I0(\rd_data[20]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[16]_i_8_n_0 ),
        .I3(\rd_data[22]_i_9_n_0 ),
        .I4(\rd_data[18]_i_8_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[16]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[16]_i_5 
       (.I0(\rd_data[16]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[20]_i_10_n_0 ),
        .I3(\rd_data[18]_i_9_n_0 ),
        .I4(\rd_data[22]_i_10_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[16]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[16]_i_6 
       (.I0(\rd_data[17]_i_10_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[16]_i_10_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [16]),
        .O(\rd_data[16]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[16]_i_7 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [16]),
        .I3(\processor/execute/alu_y [16]),
        .O(\rd_data[16]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    \rd_data[16]_i_8 
       (.I0(\processor/execute/alu_x [24]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [31]),
        .I3(\processor/execute/alu_y [4]),
        .I4(\processor/execute/alu_x [16]),
        .O(\rd_data[16]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \rd_data[16]_i_9 
       (.I0(\processor/execute/alu_x [1]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [9]),
        .I3(\processor/execute/alu_y [4]),
        .O(\rd_data[16]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[17]_i_1 
       (.I0(\rd_data[17]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[17]_i_3_n_0 ),
        .O(\processor/ex_rd_data [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[17]_i_10 
       (.I0(\rd_data[17]_i_12_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[17]_i_13_n_0 ),
        .I3(\rd_data[19]_i_23_n_0 ),
        .I4(\rd_data[19]_i_24_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[17]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[17]_i_11 
       (.I0(\rd_data[17]_i_14_n_0 ),
        .I1(\csr_data_out[17]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [17]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \rd_data[17]_i_12 
       (.I0(\processor/execute/alu_x [29]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [21]),
        .I3(\processor/execute/alu_y [4]),
        .O(\rd_data[17]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \rd_data[17]_i_13 
       (.I0(\processor/execute/alu_x [25]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [17]),
        .I3(\processor/execute/alu_y [4]),
        .O(\rd_data[17]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[17]_i_14 
       (.I0(\processor/ex_pc [17]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [17]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [17]),
        .O(\rd_data[17]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[17]_i_2 
       (.I0(\rd_data[18]_i_4_n_0 ),
        .I1(\rd_data[17]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[17]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[18]_i_5_n_0 ),
        .O(\rd_data[17]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[17]_i_3 
       (.I0(\rd_data[17]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [17]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[17]_i_7_n_0 ),
        .O(\rd_data[17]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[17]_i_4 
       (.I0(\rd_data[21]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[17]_i_8_n_0 ),
        .I3(\rd_data[19]_i_9_n_0 ),
        .I4(\rd_data[19]_i_10_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[17]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[17]_i_5 
       (.I0(\rd_data[17]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[21]_i_10_n_0 ),
        .I3(\rd_data[19]_i_11_n_0 ),
        .I4(\rd_data[23]_i_10_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[17]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[17]_i_6 
       (.I0(\rd_data[18]_i_10_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[17]_i_10_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [17]),
        .O(\rd_data[17]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[17]_i_7 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [17]),
        .I3(\processor/execute/alu_y [17]),
        .O(\rd_data[17]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    \rd_data[17]_i_8 
       (.I0(\processor/execute/alu_x [25]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [31]),
        .I3(\processor/execute/alu_y [4]),
        .I4(\processor/execute/alu_x [17]),
        .O(\rd_data[17]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \rd_data[17]_i_9 
       (.I0(\processor/execute/alu_x [2]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [10]),
        .I3(\processor/execute/alu_y [4]),
        .O(\rd_data[17]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[18]_i_1 
       (.I0(\rd_data[18]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[18]_i_3_n_0 ),
        .O(\processor/ex_rd_data [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \rd_data[18]_i_10 
       (.I0(\rd_data[18]_i_12_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[18]_i_13_n_0 ),
        .I3(\rd_data[20]_i_13_n_0 ),
        .I4(\processor/execute/alu_y [1]),
        .O(\rd_data[18]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[18]_i_11 
       (.I0(\rd_data[18]_i_14_n_0 ),
        .I1(\csr_data_out[18]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [18]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \rd_data[18]_i_12 
       (.I0(\processor/execute/alu_x [30]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [22]),
        .I3(\processor/execute/alu_y [4]),
        .O(\rd_data[18]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \rd_data[18]_i_13 
       (.I0(\processor/execute/alu_x [26]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [18]),
        .I3(\processor/execute/alu_y [4]),
        .O(\rd_data[18]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[18]_i_14 
       (.I0(\processor/ex_pc [18]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [18]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [18]),
        .O(\rd_data[18]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[18]_i_2 
       (.I0(\rd_data[19]_i_4_n_0 ),
        .I1(\rd_data[18]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[18]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[19]_i_5_n_0 ),
        .O(\rd_data[18]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[18]_i_3 
       (.I0(\rd_data[18]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [18]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[18]_i_7_n_0 ),
        .O(\rd_data[18]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[18]_i_4 
       (.I0(\rd_data[22]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[18]_i_8_n_0 ),
        .I3(\rd_data[20]_i_8_n_0 ),
        .I4(\rd_data[20]_i_9_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[18]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[18]_i_5 
       (.I0(\rd_data[18]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[22]_i_10_n_0 ),
        .I3(\rd_data[20]_i_10_n_0 ),
        .I4(\rd_data[24]_i_9_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[18]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[18]_i_6 
       (.I0(\rd_data[19]_i_12_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[18]_i_10_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [18]),
        .O(\rd_data[18]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[18]_i_7 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [18]),
        .I3(\processor/execute/alu_y [18]),
        .O(\rd_data[18]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    \rd_data[18]_i_8 
       (.I0(\processor/execute/alu_x [26]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [31]),
        .I3(\processor/execute/alu_y [4]),
        .I4(\processor/execute/alu_x [18]),
        .O(\rd_data[18]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2320)) 
    \rd_data[18]_i_9 
       (.I0(\processor/execute/alu_x [3]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_x [11]),
        .O(\rd_data[18]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[19]_i_1 
       (.I0(\rd_data[19]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[19]_i_3_n_0 ),
        .O(\processor/ex_rd_data [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    \rd_data[19]_i_10 
       (.I0(\processor/execute/alu_x [27]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [31]),
        .I3(\processor/execute/alu_y [4]),
        .I4(\processor/execute/alu_x [19]),
        .O(\rd_data[19]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \rd_data[19]_i_11 
       (.I0(\processor/execute/alu_x [4]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [12]),
        .I3(\processor/execute/alu_y [4]),
        .O(\rd_data[19]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \rd_data[19]_i_12 
       (.I0(\rd_data[19]_i_23_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[19]_i_24_n_0 ),
        .I3(\rd_data[21]_i_13_n_0 ),
        .I4(\processor/execute/alu_y [1]),
        .O(\rd_data[19]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[19]_i_14 
       (.I0(\rd_data[19]_i_29_n_0 ),
        .I1(\rd_data[19]_i_30_n_0 ),
        .I2(\rd_data[19]_i_31_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [19]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[19]_i_15 
       (.I0(\rd_data[19]_i_32_n_0 ),
        .I1(\rd_data[19]_i_33_n_0 ),
        .I2(\rd_data[19]_i_34_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [18]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[19]_i_16 
       (.I0(\rd_data[19]_i_35_n_0 ),
        .I1(\rd_data[19]_i_36_n_0 ),
        .I2(\rd_data[19]_i_37_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [17]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[19]_i_17 
       (.I0(\rd_data[19]_i_38_n_0 ),
        .I1(\rd_data[19]_i_39_n_0 ),
        .I2(\rd_data[19]_i_40_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [16]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[19]_i_18 
       (.I0(\processor/execute/alu_x [19]),
        .I1(\processor/execute/alu_y [19]),
        .O(\rd_data[19]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[19]_i_19 
       (.I0(\processor/execute/alu_x [18]),
        .I1(\processor/execute/alu_y [18]),
        .O(\rd_data[19]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[19]_i_2 
       (.I0(\rd_data[20]_i_4_n_0 ),
        .I1(\rd_data[19]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[19]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[20]_i_5_n_0 ),
        .O(\rd_data[19]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[19]_i_20 
       (.I0(\processor/execute/alu_x [17]),
        .I1(\processor/execute/alu_y [17]),
        .O(\rd_data[19]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[19]_i_21 
       (.I0(\processor/execute/alu_x [16]),
        .I1(\processor/execute/alu_y [16]),
        .O(\rd_data[19]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[19]_i_22 
       (.I0(\rd_data[19]_i_42_n_0 ),
        .I1(\csr_data_out[19]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [19]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \rd_data[19]_i_23 
       (.I0(\processor/execute/alu_x [31]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [23]),
        .I3(\processor/execute/alu_y [4]),
        .O(\rd_data[19]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \rd_data[19]_i_24 
       (.I0(\processor/execute/alu_x [27]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [19]),
        .I3(\processor/execute/alu_y [4]),
        .O(\rd_data[19]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[19]_i_25 
       (.I0(\processor/execute/alu_x [19]),
        .I1(\processor/execute/alu_y [19]),
        .O(\rd_data[19]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[19]_i_26 
       (.I0(\processor/execute/alu_x [18]),
        .I1(\processor/execute/alu_y [18]),
        .O(\rd_data[19]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[19]_i_27 
       (.I0(\processor/execute/alu_x [17]),
        .I1(\processor/execute/alu_y [17]),
        .O(\rd_data[19]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[19]_i_28 
       (.I0(\processor/execute/alu_x [16]),
        .I1(\processor/execute/alu_y [16]),
        .O(\rd_data[19]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[19]_i_29 
       (.I0(\processor/ex_pc [19]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [19]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [19]),
        .O(\rd_data[19]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[19]_i_3 
       (.I0(\rd_data[19]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [19]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[19]_i_8_n_0 ),
        .O(\rd_data[19]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rd_data[19]_i_30 
       (.I0(\processor/mem_exception_context[badaddr] [19]),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .O(\rd_data[19]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000540455555555)) 
    \rd_data[19]_i_31 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\rd_data[19]_i_43_n_0 ),
        .I2(\csr_data_out[30]_i_9_n_0 ),
        .I3(\processor/wb_exception_context[badaddr] [19]),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\rd_data[19]_i_44_n_0 ),
        .O(\rd_data[19]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[19]_i_32 
       (.I0(\processor/ex_pc [18]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [18]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [18]),
        .O(\rd_data[19]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rd_data[19]_i_33 
       (.I0(\processor/mem_exception_context[badaddr] [18]),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .O(\rd_data[19]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000540455555555)) 
    \rd_data[19]_i_34 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\rd_data[19]_i_45_n_0 ),
        .I2(\csr_data_out[30]_i_9_n_0 ),
        .I3(\processor/wb_exception_context[badaddr] [18]),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\rd_data[19]_i_46_n_0 ),
        .O(\rd_data[19]_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[19]_i_35 
       (.I0(\processor/ex_pc [17]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [17]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [17]),
        .O(\rd_data[19]_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rd_data[19]_i_36 
       (.I0(\processor/mem_exception_context[badaddr] [17]),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .O(\rd_data[19]_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000540455555555)) 
    \rd_data[19]_i_37 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\rd_data[19]_i_47_n_0 ),
        .I2(\csr_data_out[30]_i_9_n_0 ),
        .I3(\processor/wb_exception_context[badaddr] [17]),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\rd_data[19]_i_48_n_0 ),
        .O(\rd_data[19]_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[19]_i_38 
       (.I0(\processor/ex_pc [16]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [16]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [16]),
        .O(\rd_data[19]_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rd_data[19]_i_39 
       (.I0(\processor/mem_exception_context[badaddr] [16]),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .O(\rd_data[19]_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[19]_i_4 
       (.I0(\rd_data[21]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[21]_i_9_n_0 ),
        .I3(\rd_data[19]_i_9_n_0 ),
        .I4(\rd_data[19]_i_10_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[19]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000540455555555)) 
    \rd_data[19]_i_40 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\rd_data[19]_i_49_n_0 ),
        .I2(\csr_data_out[30]_i_9_n_0 ),
        .I3(\processor/wb_exception_context[badaddr] [16]),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\rd_data[19]_i_50_n_0 ),
        .O(\rd_data[19]_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[19]_i_42 
       (.I0(\processor/ex_pc [19]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [19]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [19]),
        .O(\rd_data[19]_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCAAACAAACAAAAAAA)) 
    \rd_data[19]_i_43 
       (.I0(\processor/csr_read_data [19]),
        .I1(\processor/wb_csr_data [19]),
        .I2(\processor/execute/csr_writeable ),
        .I3(\processor/execute/csr_value_forwarded3 ),
        .I4(\processor/wb_csr_write [1]),
        .I5(\processor/wb_csr_write [0]),
        .O(\rd_data[19]_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7F7F7FFF)) 
    \rd_data[19]_i_44 
       (.I0(\processor/mem_csr_data [19]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/mem_csr_write [0]),
        .I4(\processor/mem_csr_write [1]),
        .O(\rd_data[19]_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCAAACAAACAAAAAAA)) 
    \rd_data[19]_i_45 
       (.I0(\processor/csr_read_data [18]),
        .I1(\processor/wb_csr_data [18]),
        .I2(\processor/execute/csr_writeable ),
        .I3(\processor/execute/csr_value_forwarded3 ),
        .I4(\processor/wb_csr_write [1]),
        .I5(\processor/wb_csr_write [0]),
        .O(\rd_data[19]_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7F7F7FFF)) 
    \rd_data[19]_i_46 
       (.I0(\processor/mem_csr_data [18]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/mem_csr_write [0]),
        .I4(\processor/mem_csr_write [1]),
        .O(\rd_data[19]_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCAAACAAACAAAAAAA)) 
    \rd_data[19]_i_47 
       (.I0(\processor/csr_read_data [17]),
        .I1(\processor/wb_csr_data [17]),
        .I2(\processor/execute/csr_writeable ),
        .I3(\processor/execute/csr_value_forwarded3 ),
        .I4(\processor/wb_csr_write [1]),
        .I5(\processor/wb_csr_write [0]),
        .O(\rd_data[19]_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7F7F7FFF)) 
    \rd_data[19]_i_48 
       (.I0(\processor/mem_csr_data [17]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/mem_csr_write [0]),
        .I4(\processor/mem_csr_write [1]),
        .O(\rd_data[19]_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCAAACAAACAAAAAAA)) 
    \rd_data[19]_i_49 
       (.I0(\processor/csr_read_data [16]),
        .I1(\processor/wb_csr_data [16]),
        .I2(\processor/execute/csr_writeable ),
        .I3(\processor/execute/csr_value_forwarded3 ),
        .I4(\processor/wb_csr_write [1]),
        .I5(\processor/wb_csr_write [0]),
        .O(\rd_data[19]_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[19]_i_5 
       (.I0(\rd_data[21]_i_10_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[25]_i_9_n_0 ),
        .I3(\rd_data[19]_i_11_n_0 ),
        .I4(\rd_data[23]_i_10_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[19]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7F7F7FFF)) 
    \rd_data[19]_i_50 
       (.I0(\processor/mem_csr_data [16]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/mem_csr_write [0]),
        .I4(\processor/mem_csr_write [1]),
        .O(\rd_data[19]_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[19]_i_6 
       (.I0(\rd_data[20]_i_11_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[19]_i_12_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [19]),
        .O(\rd_data[19]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[19]_i_8 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [19]),
        .I3(\processor/execute/alu_y [19]),
        .O(\rd_data[19]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hCDC8)) 
    \rd_data[19]_i_9 
       (.I0(\processor/execute/alu_y [3]),
        .I1(\processor/execute/alu_x [31]),
        .I2(\processor/execute/alu_y [4]),
        .I3(\processor/execute/alu_x [23]),
        .O(\rd_data[19]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[1]_i_10 
       (.I0(\processor/execute/alu_x [26]),
        .I1(\processor/execute/alu_x [10]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_x [18]),
        .I4(\processor/execute/alu_y [4]),
        .I5(\processor/execute/alu_x [2]),
        .O(\rd_data[1]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[1]_i_11 
       (.I0(\processor/execute/alu_x [27]),
        .I1(\processor/execute/alu_x [11]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_x [19]),
        .I4(\processor/execute/alu_y [4]),
        .I5(\processor/execute/alu_x [3]),
        .O(\rd_data[1]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[1]_i_12 
       (.I0(\processor/execute/alu_x [25]),
        .I1(\processor/execute/alu_x [9]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_x [17]),
        .I4(\processor/execute/alu_y [4]),
        .I5(\processor/execute/alu_x [1]),
        .O(\rd_data[1]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[1]_i_2 
       (.I0(\rd_data[1]_i_4_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [1]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[1]_i_5_n_0 ),
        .O(\rd_data[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \rd_data[1]_i_3 
       (.I0(\rd_data[2]_i_7_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[1]_i_6_n_0 ),
        .I3(\rd_data[31]_i_10_n_0 ),
        .I4(\processor/execute/alu_instance/data9 [1]),
        .I5(\rd_data[31]_i_11_n_0 ),
        .O(\rd_data[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[1]_i_4 
       (.I0(\rd_data[1]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[1]_i_9_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [1]),
        .O(\rd_data[1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[1]_i_5 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [1]),
        .I3(\processor/execute/alu_y [1]),
        .O(\rd_data[1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000002)) 
    \rd_data[1]_i_6 
       (.I0(\processor/execute/alu_x [0]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_y [2]),
        .I3(\processor/execute/alu_y [3]),
        .I4(\processor/execute/alu_y [1]),
        .O(\rd_data[1]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[1]_i_7 
       (.I0(\rd_data[4]_i_8_n_0_repN ),
        .I1(\processor/execute/alu_y [1]),
        .I2(\rd_data[2]_i_14_n_0 ),
        .I3(\processor/execute/alu_y [0]),
        .I4(\rd_data[1]_i_9_n_0 ),
        .O(\processor/execute/alu_instance/data9 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[1]_i_8 
       (.I0(\rd_data[8]_i_12_n_0 ),
        .I1(\rd_data[4]_i_11_n_0 ),
        .I2(\processor/execute/alu_y [1]),
        .I3(\rd_data[6]_i_8_n_0 ),
        .I4(\processor/execute/alu_y [2]),
        .I5(\rd_data[1]_i_10_n_0 ),
        .O(\rd_data[1]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[1]_i_9 
       (.I0(\rd_data[7]_i_9_n_0 ),
        .I1(\rd_data[1]_i_11_n_0 ),
        .I2(\processor/execute/alu_y [1]),
        .I3(\rd_data[5]_i_8_n_0 ),
        .I4(\processor/execute/alu_y [2]),
        .I5(\rd_data[1]_i_12_n_0 ),
        .O(\rd_data[1]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[20]_i_1 
       (.I0(\rd_data[20]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[20]_i_3_n_0 ),
        .O(\processor/ex_rd_data [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \rd_data[20]_i_10 
       (.I0(\processor/execute/alu_x [5]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [13]),
        .I3(\processor/execute/alu_y [4]),
        .O(\rd_data[20]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rd_data[20]_i_11 
       (.I0(\rd_data[22]_i_13_n_0 ),
        .I1(\processor/execute/alu_y [1]),
        .I2(\rd_data[20]_i_13_n_0 ),
        .O(\rd_data[20]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[20]_i_12 
       (.I0(\rd_data[20]_i_14_n_0 ),
        .I1(\csr_data_out[20]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [20]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h04FF0400)) 
    \rd_data[20]_i_13 
       (.I0(\processor/execute/alu_y [4]),
        .I1(\processor/execute/alu_x [24]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_y [2]),
        .I4(\rd_data[16]_i_12_n_0 ),
        .O(\rd_data[20]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[20]_i_14 
       (.I0(\processor/ex_pc [20]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [20]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [20]),
        .O(\rd_data[20]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[20]_i_2 
       (.I0(\rd_data[21]_i_4_n_0 ),
        .I1(\rd_data[20]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[20]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[21]_i_5_n_0 ),
        .O(\rd_data[20]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[20]_i_3 
       (.I0(\rd_data[20]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [20]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[20]_i_7_n_0 ),
        .O(\rd_data[20]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[20]_i_4 
       (.I0(\rd_data[22]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[22]_i_9_n_0 ),
        .I3(\rd_data[20]_i_8_n_0 ),
        .I4(\rd_data[20]_i_9_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[20]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[20]_i_5 
       (.I0(\rd_data[20]_i_10_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[24]_i_9_n_0 ),
        .I3(\rd_data[22]_i_10_n_0 ),
        .I4(\rd_data[26]_i_9_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[20]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[20]_i_6 
       (.I0(\rd_data[21]_i_11_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[20]_i_11_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [20]),
        .O(\rd_data[20]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[20]_i_7 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [20]),
        .I3(\processor/execute/alu_y [20]),
        .O(\rd_data[20]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hCDC8)) 
    \rd_data[20]_i_8 
       (.I0(\processor/execute/alu_y [3]),
        .I1(\processor/execute/alu_x [31]),
        .I2(\processor/execute/alu_y [4]),
        .I3(\processor/execute/alu_x [24]),
        .O(\rd_data[20]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    \rd_data[20]_i_9 
       (.I0(\processor/execute/alu_x [28]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [31]),
        .I3(\processor/execute/alu_y [4]),
        .I4(\processor/execute/alu_x [20]),
        .O(\rd_data[20]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[21]_i_1 
       (.I0(\rd_data[21]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[21]_i_3_n_0 ),
        .O(\processor/ex_rd_data [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \rd_data[21]_i_10 
       (.I0(\processor/execute/alu_x [6]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [14]),
        .I3(\processor/execute/alu_y [4]),
        .O(\rd_data[21]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rd_data[21]_i_11 
       (.I0(\rd_data[23]_i_22_n_0 ),
        .I1(\processor/execute/alu_y [1]),
        .I2(\rd_data[21]_i_13_n_0 ),
        .O(\rd_data[21]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[21]_i_12 
       (.I0(\rd_data[21]_i_14_n_0 ),
        .I1(\csr_data_out[21]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [21]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h04FF0400)) 
    \rd_data[21]_i_13 
       (.I0(\processor/execute/alu_y [4]),
        .I1(\processor/execute/alu_x [25]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_y [2]),
        .I4(\rd_data[17]_i_12_n_0 ),
        .O(\rd_data[21]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[21]_i_14 
       (.I0(\processor/ex_pc [21]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [21]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [21]),
        .O(\rd_data[21]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[21]_i_2 
       (.I0(\rd_data[22]_i_4_n_0 ),
        .I1(\rd_data[21]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[21]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[22]_i_5_n_0 ),
        .O(\rd_data[21]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[21]_i_3 
       (.I0(\rd_data[21]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [21]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[21]_i_7_n_0 ),
        .O(\rd_data[21]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \rd_data[21]_i_4 
       (.I0(\rd_data[21]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[21]_i_9_n_0 ),
        .I3(\rd_data[23]_i_9_n_0 ),
        .I4(\processor/execute/alu_y [1]),
        .O(\rd_data[21]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[21]_i_5 
       (.I0(\rd_data[21]_i_10_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[25]_i_9_n_0 ),
        .I3(\rd_data[23]_i_10_n_0 ),
        .I4(\rd_data[27]_i_11_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[21]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[21]_i_6 
       (.I0(\rd_data[22]_i_11_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[21]_i_11_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [21]),
        .O(\rd_data[21]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[21]_i_7 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [21]),
        .I3(\processor/execute/alu_y [21]),
        .O(\rd_data[21]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hCDC8)) 
    \rd_data[21]_i_8 
       (.I0(\processor/execute/alu_y [3]),
        .I1(\processor/execute/alu_x [31]),
        .I2(\processor/execute/alu_y [4]),
        .I3(\processor/execute/alu_x [25]),
        .O(\rd_data[21]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    \rd_data[21]_i_9 
       (.I0(\processor/execute/alu_x [29]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [31]),
        .I3(\processor/execute/alu_y [4]),
        .I4(\processor/execute/alu_x [21]),
        .O(\rd_data[21]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[22]_i_1 
       (.I0(\rd_data[22]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[22]_i_3_n_0 ),
        .O(\processor/ex_rd_data [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \rd_data[22]_i_10 
       (.I0(\processor/execute/alu_x [7]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [15]),
        .I3(\processor/execute/alu_y [4]),
        .O(\rd_data[22]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rd_data[22]_i_11 
       (.I0(\rd_data[24]_i_12_n_0 ),
        .I1(\processor/execute/alu_y [1]),
        .I2(\rd_data[22]_i_13_n_0 ),
        .O(\rd_data[22]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[22]_i_12 
       (.I0(\rd_data[22]_i_14_n_0 ),
        .I1(\csr_data_out[22]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [22]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h04FF0400)) 
    \rd_data[22]_i_13 
       (.I0(\processor/execute/alu_y [4]),
        .I1(\processor/execute/alu_x [26]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_y [2]),
        .I4(\rd_data[18]_i_12_n_0 ),
        .O(\rd_data[22]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[22]_i_14 
       (.I0(\processor/ex_pc [22]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [22]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [22]),
        .O(\rd_data[22]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[22]_i_2 
       (.I0(\rd_data[23]_i_4_n_0 ),
        .I1(\rd_data[22]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[22]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[23]_i_5_n_0 ),
        .O(\rd_data[22]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[22]_i_3 
       (.I0(\rd_data[22]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [22]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[22]_i_7_n_0 ),
        .O(\rd_data[22]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \rd_data[22]_i_4 
       (.I0(\rd_data[22]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[22]_i_9_n_0 ),
        .I3(\rd_data[24]_i_8_n_0 ),
        .I4(\processor/execute/alu_y [1]),
        .O(\rd_data[22]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[22]_i_5 
       (.I0(\rd_data[22]_i_10_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[26]_i_9_n_0 ),
        .I3(\rd_data[24]_i_9_n_0 ),
        .I4(\rd_data[28]_i_10_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[22]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[22]_i_6 
       (.I0(\rd_data[23]_i_11_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[22]_i_11_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [22]),
        .O(\rd_data[22]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[22]_i_7 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [22]),
        .I3(\processor/execute/alu_y [22]),
        .O(\rd_data[22]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hCDC8)) 
    \rd_data[22]_i_8 
       (.I0(\processor/execute/alu_y [3]),
        .I1(\processor/execute/alu_x [31]),
        .I2(\processor/execute/alu_y [4]),
        .I3(\processor/execute/alu_x [26]),
        .O(\rd_data[22]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    \rd_data[22]_i_9 
       (.I0(\processor/execute/alu_x [30]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [31]),
        .I3(\processor/execute/alu_y [4]),
        .I4(\processor/execute/alu_x [22]),
        .O(\rd_data[22]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[23]_i_1 
       (.I0(\rd_data[23]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[23]_i_3_n_0 ),
        .O(\processor/ex_rd_data [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h3300B8B8)) 
    \rd_data[23]_i_10 
       (.I0(\processor/execute/alu_x [0]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [16]),
        .I3(\processor/execute/alu_x [8]),
        .I4(\processor/execute/alu_y [3]),
        .O(\rd_data[23]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rd_data[23]_i_11 
       (.I0(\rd_data[25]_i_12_n_0 ),
        .I1(\processor/execute/alu_y [1]),
        .I2(\rd_data[23]_i_22_n_0 ),
        .O(\rd_data[23]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[23]_i_13 
       (.I0(\rd_data[23]_i_27_n_0 ),
        .I1(\rd_data[23]_i_28_n_0 ),
        .I2(\rd_data[23]_i_29_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [23]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[23]_i_14 
       (.I0(\rd_data[23]_i_30_n_0 ),
        .I1(\rd_data[23]_i_31_n_0 ),
        .I2(\rd_data[23]_i_32_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [22]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[23]_i_15 
       (.I0(\rd_data[23]_i_33_n_0 ),
        .I1(\rd_data[23]_i_34_n_0 ),
        .I2(\rd_data[23]_i_35_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [21]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[23]_i_16 
       (.I0(\rd_data[23]_i_36_n_0 ),
        .I1(\rd_data[23]_i_37_n_0 ),
        .I2(\rd_data[23]_i_38_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [20]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[23]_i_17 
       (.I0(\processor/execute/alu_x [23]),
        .I1(\processor/execute/alu_y [23]),
        .O(\rd_data[23]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[23]_i_18 
       (.I0(\processor/execute/alu_x [22]),
        .I1(\processor/execute/alu_y [22]),
        .O(\rd_data[23]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[23]_i_19 
       (.I0(\processor/execute/alu_x [21]),
        .I1(\processor/execute/alu_y [21]),
        .O(\rd_data[23]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[23]_i_2 
       (.I0(\rd_data[24]_i_4_n_0 ),
        .I1(\rd_data[23]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[23]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[24]_i_5_n_0 ),
        .O(\rd_data[23]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[23]_i_20 
       (.I0(\processor/execute/alu_x [20]),
        .I1(\processor/execute/alu_y [20]),
        .O(\rd_data[23]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[23]_i_21 
       (.I0(\rd_data[23]_i_40_n_0 ),
        .I1(\csr_data_out[23]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [23]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \rd_data[23]_i_22 
       (.I0(\processor/execute/alu_x [27]),
        .I1(\processor/execute/alu_y [2]),
        .I2(\processor/execute/alu_x [31]),
        .I3(\processor/execute/alu_y [3]),
        .I4(\processor/execute/alu_x [23]),
        .I5(\processor/execute/alu_y [4]),
        .O(\rd_data[23]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[23]_i_23 
       (.I0(\processor/execute/alu_x [23]),
        .I1(\processor/execute/alu_y [23]),
        .O(\rd_data[23]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[23]_i_24 
       (.I0(\processor/execute/alu_x [22]),
        .I1(\processor/execute/alu_y [22]),
        .O(\rd_data[23]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[23]_i_25 
       (.I0(\processor/execute/alu_x [21]),
        .I1(\processor/execute/alu_y [21]),
        .O(\rd_data[23]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[23]_i_26 
       (.I0(\processor/execute/alu_x [20]),
        .I1(\processor/execute/alu_y [20]),
        .O(\rd_data[23]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[23]_i_27 
       (.I0(\processor/ex_pc [23]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [23]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [23]),
        .O(\rd_data[23]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rd_data[23]_i_28 
       (.I0(\processor/mem_exception_context[badaddr] [23]),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .O(\rd_data[23]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000540455555555)) 
    \rd_data[23]_i_29 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\rd_data[23]_i_41_n_0 ),
        .I2(\csr_data_out[30]_i_9_n_0 ),
        .I3(\processor/wb_exception_context[badaddr] [23]),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\rd_data[23]_i_42_n_0 ),
        .O(\rd_data[23]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[23]_i_3 
       (.I0(\rd_data[23]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [23]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[23]_i_8_n_0 ),
        .O(\rd_data[23]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[23]_i_30 
       (.I0(\processor/ex_pc [22]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [22]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [22]),
        .O(\rd_data[23]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rd_data[23]_i_31 
       (.I0(\processor/mem_exception_context[badaddr] [22]),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .O(\rd_data[23]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000540455555555)) 
    \rd_data[23]_i_32 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\rd_data[23]_i_43_n_0 ),
        .I2(\csr_data_out[30]_i_9_n_0 ),
        .I3(\processor/wb_exception_context[badaddr] [22]),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\rd_data[23]_i_44_n_0 ),
        .O(\rd_data[23]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[23]_i_33 
       (.I0(\processor/ex_pc [21]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [21]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [21]),
        .O(\rd_data[23]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rd_data[23]_i_34 
       (.I0(\processor/mem_exception_context[badaddr] [21]),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .O(\rd_data[23]_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000540455555555)) 
    \rd_data[23]_i_35 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\rd_data[23]_i_45_n_0 ),
        .I2(\csr_data_out[30]_i_9_n_0 ),
        .I3(\processor/wb_exception_context[badaddr] [21]),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\rd_data[23]_i_46_n_0 ),
        .O(\rd_data[23]_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[23]_i_36 
       (.I0(\processor/ex_pc [20]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [20]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [20]),
        .O(\rd_data[23]_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rd_data[23]_i_37 
       (.I0(\processor/mem_exception_context[badaddr] [20]),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .O(\rd_data[23]_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000540455555555)) 
    \rd_data[23]_i_38 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\rd_data[23]_i_47_n_0 ),
        .I2(\csr_data_out[30]_i_9_n_0 ),
        .I3(\processor/wb_exception_context[badaddr] [20]),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\rd_data[23]_i_48_n_0 ),
        .O(\rd_data[23]_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rd_data[23]_i_4 
       (.I0(\rd_data[25]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [1]),
        .I2(\rd_data[23]_i_9_n_0 ),
        .O(\rd_data[23]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[23]_i_40 
       (.I0(\processor/ex_pc [23]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [23]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [23]),
        .O(\rd_data[23]_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCAAACAAACAAAAAAA)) 
    \rd_data[23]_i_41 
       (.I0(\processor/csr_read_data [23]),
        .I1(\processor/wb_csr_data [23]),
        .I2(\processor/execute/csr_writeable ),
        .I3(\processor/execute/csr_value_forwarded3 ),
        .I4(\processor/wb_csr_write [1]),
        .I5(\processor/wb_csr_write [0]),
        .O(\rd_data[23]_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7F7F7FFF)) 
    \rd_data[23]_i_42 
       (.I0(\processor/mem_csr_data [23]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/mem_csr_write [0]),
        .I4(\processor/mem_csr_write [1]),
        .O(\rd_data[23]_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCAAACAAACAAAAAAA)) 
    \rd_data[23]_i_43 
       (.I0(\processor/csr_read_data [22]),
        .I1(\processor/wb_csr_data [22]),
        .I2(\processor/execute/csr_writeable ),
        .I3(\processor/execute/csr_value_forwarded3 ),
        .I4(\processor/wb_csr_write [1]),
        .I5(\processor/wb_csr_write [0]),
        .O(\rd_data[23]_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7F7F7FFF)) 
    \rd_data[23]_i_44 
       (.I0(\processor/mem_csr_data [22]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/mem_csr_write [0]),
        .I4(\processor/mem_csr_write [1]),
        .O(\rd_data[23]_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCAAACAAACAAAAAAA)) 
    \rd_data[23]_i_45 
       (.I0(\processor/csr_read_data [21]),
        .I1(\processor/wb_csr_data [21]),
        .I2(\processor/execute/csr_writeable ),
        .I3(\processor/execute/csr_value_forwarded3 ),
        .I4(\processor/wb_csr_write [1]),
        .I5(\processor/wb_csr_write [0]),
        .O(\rd_data[23]_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7F7F7FFF)) 
    \rd_data[23]_i_46 
       (.I0(\processor/mem_csr_data [21]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/mem_csr_write [0]),
        .I4(\processor/mem_csr_write [1]),
        .O(\rd_data[23]_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCAAACAAACAAAAAAA)) 
    \rd_data[23]_i_47 
       (.I0(\processor/csr_read_data [20]),
        .I1(\processor/wb_csr_data [20]),
        .I2(\processor/execute/csr_writeable ),
        .I3(\processor/execute/csr_value_forwarded3 ),
        .I4(\processor/wb_csr_write [1]),
        .I5(\processor/wb_csr_write [0]),
        .O(\rd_data[23]_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7F7F7FFF)) 
    \rd_data[23]_i_48 
       (.I0(\processor/mem_csr_data [20]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/mem_csr_write [0]),
        .I4(\processor/mem_csr_write [1]),
        .O(\rd_data[23]_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[23]_i_5 
       (.I0(\rd_data[25]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[29]_i_8_n_0 ),
        .I3(\rd_data[23]_i_10_n_0 ),
        .I4(\rd_data[27]_i_11_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[23]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[23]_i_6 
       (.I0(\rd_data[24]_i_10_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[23]_i_11_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [23]),
        .O(\rd_data[23]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[23]_i_8 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [23]),
        .I3(\processor/execute/alu_y [23]),
        .O(\rd_data[23]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00FB0BFF00F808)) 
    \rd_data[23]_i_9 
       (.I0(\processor/execute/alu_x [27]),
        .I1(\processor/execute/alu_y [2]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_x [31]),
        .I4(\processor/execute/alu_y [4]),
        .I5(\processor/execute/alu_x [23]),
        .O(\rd_data[23]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[24]_i_1 
       (.I0(\rd_data[24]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[24]_i_3_n_0 ),
        .O(\processor/ex_rd_data [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rd_data[24]_i_10 
       (.I0(\rd_data[26]_i_12_n_0 ),
        .I1(\processor/execute/alu_y [1]),
        .I2(\rd_data[24]_i_12_n_0 ),
        .O(\rd_data[24]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[24]_i_11 
       (.I0(\rd_data[24]_i_13_n_0 ),
        .I1(\csr_data_out[24]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [24]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \rd_data[24]_i_12 
       (.I0(\processor/execute/alu_x [28]),
        .I1(\processor/execute/alu_y [2]),
        .I2(\processor/execute/alu_y [4]),
        .I3(\processor/execute/alu_x [24]),
        .I4(\processor/execute/alu_y [3]),
        .O(\rd_data[24]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[24]_i_13 
       (.I0(\processor/ex_pc [24]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [24]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [24]),
        .O(\rd_data[24]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[24]_i_2 
       (.I0(\rd_data[25]_i_4_n_0 ),
        .I1(\rd_data[24]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[24]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[25]_i_5_n_0 ),
        .O(\rd_data[24]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[24]_i_3 
       (.I0(\rd_data[24]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [24]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[24]_i_7_n_0 ),
        .O(\rd_data[24]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rd_data[24]_i_4 
       (.I0(\rd_data[26]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [1]),
        .I2(\rd_data[24]_i_8_n_0 ),
        .O(\rd_data[24]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[24]_i_5 
       (.I0(\rd_data[24]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[28]_i_10_n_0 ),
        .I3(\rd_data[26]_i_9_n_0 ),
        .I4(\rd_data[30]_i_12_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[24]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[24]_i_6 
       (.I0(\rd_data[25]_i_10_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[24]_i_10_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [24]),
        .O(\rd_data[24]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[24]_i_7 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [24]),
        .I3(\processor/execute/alu_y [24]),
        .O(\rd_data[24]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00FB0BFF00F808)) 
    \rd_data[24]_i_8 
       (.I0(\processor/execute/alu_x [28]),
        .I1(\processor/execute/alu_y [2]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_x [31]),
        .I4(\processor/execute/alu_y [4]),
        .I5(\processor/execute/alu_x [24]),
        .O(\rd_data[24]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h3300B8B8)) 
    \rd_data[24]_i_9 
       (.I0(\processor/execute/alu_x [1]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [17]),
        .I3(\processor/execute/alu_x [9]),
        .I4(\processor/execute/alu_y [3]),
        .O(\rd_data[24]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[25]_i_1 
       (.I0(\rd_data[25]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[25]_i_3_n_0 ),
        .O(\processor/ex_rd_data [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rd_data[25]_i_10 
       (.I0(\rd_data[27]_i_23_n_0 ),
        .I1(\processor/execute/alu_y [1]),
        .I2(\rd_data[25]_i_12_n_0 ),
        .O(\rd_data[25]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[25]_i_11 
       (.I0(\rd_data[25]_i_13_n_0 ),
        .I1(\csr_data_out[25]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [25]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \rd_data[25]_i_12 
       (.I0(\processor/execute/alu_x [29]),
        .I1(\processor/execute/alu_y [2]),
        .I2(\processor/execute/alu_y [4]),
        .I3(\processor/execute/alu_x [25]),
        .I4(\processor/execute/alu_y [3]),
        .O(\rd_data[25]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[25]_i_13 
       (.I0(\processor/ex_pc [25]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [25]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [25]),
        .O(\rd_data[25]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[25]_i_2 
       (.I0(\rd_data[26]_i_4_n_0 ),
        .I1(\rd_data[25]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[25]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[26]_i_5_n_0 ),
        .O(\rd_data[25]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[25]_i_3 
       (.I0(\rd_data[25]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [25]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[25]_i_7_n_0 ),
        .O(\rd_data[25]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rd_data[25]_i_4 
       (.I0(\rd_data[27]_i_10_n_0 ),
        .I1(\processor/execute/alu_y [1]),
        .I2(\rd_data[25]_i_8_n_0 ),
        .O(\rd_data[25]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[25]_i_5 
       (.I0(\rd_data[25]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[29]_i_8_n_0 ),
        .I3(\rd_data[27]_i_11_n_0 ),
        .I4(\rd_data[31]_i_24_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[25]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[25]_i_6 
       (.I0(\rd_data[26]_i_10_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[25]_i_10_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [25]),
        .O(\rd_data[25]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[25]_i_7 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [25]),
        .I3(\processor/execute/alu_y [25]),
        .O(\rd_data[25]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00FB0BFF00F808)) 
    \rd_data[25]_i_8 
       (.I0(\processor/execute/alu_x [29]),
        .I1(\processor/execute/alu_y [2]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_x [31]),
        .I4(\processor/execute/alu_y [4]),
        .I5(\processor/execute/alu_x [25]),
        .O(\rd_data[25]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h3300B8B8)) 
    \rd_data[25]_i_9 
       (.I0(\processor/execute/alu_x [2]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [18]),
        .I3(\processor/execute/alu_x [10]),
        .I4(\processor/execute/alu_y [3]),
        .O(\rd_data[25]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[26]_i_1 
       (.I0(\rd_data[26]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[26]_i_3_n_0 ),
        .O(\processor/ex_rd_data [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \rd_data[26]_i_10 
       (.I0(\processor/execute/alu_y [3]),
        .I1(\processor/execute/alu_x [28]),
        .I2(\processor/execute/alu_y [4]),
        .I3(\processor/execute/alu_y [2]),
        .I4(\processor/execute/alu_y [1]),
        .I5(\rd_data[26]_i_12_n_0 ),
        .O(\rd_data[26]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[26]_i_11 
       (.I0(\rd_data[26]_i_13_n_0 ),
        .I1(\csr_data_out[26]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [26]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \rd_data[26]_i_12 
       (.I0(\processor/execute/alu_x [30]),
        .I1(\processor/execute/alu_y [2]),
        .I2(\processor/execute/alu_y [4]),
        .I3(\processor/execute/alu_x [26]),
        .I4(\processor/execute/alu_y [3]),
        .O(\rd_data[26]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[26]_i_13 
       (.I0(\processor/ex_pc [26]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [26]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [26]),
        .O(\rd_data[26]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[26]_i_2 
       (.I0(\rd_data[27]_i_4_n_0 ),
        .I1(\rd_data[26]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[26]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[27]_i_5_n_0 ),
        .O(\rd_data[26]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[26]_i_3 
       (.I0(\rd_data[26]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [26]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[26]_i_7_n_0 ),
        .O(\rd_data[26]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rd_data[26]_i_4 
       (.I0(\rd_data[28]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [1]),
        .I2(\rd_data[26]_i_8_n_0 ),
        .O(\rd_data[26]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[26]_i_5 
       (.I0(\rd_data[26]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[30]_i_12_n_0 ),
        .I3(\rd_data[28]_i_10_n_0 ),
        .I4(\rd_data[31]_i_18_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[26]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[26]_i_6 
       (.I0(\rd_data[27]_i_12_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[26]_i_10_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [26]),
        .O(\rd_data[26]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[26]_i_7 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [26]),
        .I3(\processor/execute/alu_y [26]),
        .O(\rd_data[26]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00FB0BFF00F808)) 
    \rd_data[26]_i_8 
       (.I0(\processor/execute/alu_x [30]),
        .I1(\processor/execute/alu_y [2]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_x [31]),
        .I4(\processor/execute/alu_y [4]),
        .I5(\processor/execute/alu_x [26]),
        .O(\rd_data[26]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h3300B8B8)) 
    \rd_data[26]_i_9 
       (.I0(\processor/execute/alu_x [3]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [19]),
        .I3(\processor/execute/alu_x [11]),
        .I4(\processor/execute/alu_y [3]),
        .O(\rd_data[26]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[27]_i_1 
       (.I0(\rd_data[27]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[27]_i_3_n_0 ),
        .O(\processor/ex_rd_data [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF0F1F0E0)) 
    \rd_data[27]_i_10 
       (.I0(\processor/execute/alu_y [2]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [31]),
        .I3(\processor/execute/alu_y [4]),
        .I4(\processor/execute/alu_x [27]),
        .O(\rd_data[27]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h3300B8B8)) 
    \rd_data[27]_i_11 
       (.I0(\processor/execute/alu_x [4]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [20]),
        .I3(\processor/execute/alu_x [12]),
        .I4(\processor/execute/alu_y [3]),
        .O(\rd_data[27]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \rd_data[27]_i_12 
       (.I0(\processor/execute/alu_y [3]),
        .I1(\processor/execute/alu_x [29]),
        .I2(\processor/execute/alu_y [4]),
        .I3(\processor/execute/alu_y [2]),
        .I4(\processor/execute/alu_y [1]),
        .I5(\rd_data[27]_i_23_n_0 ),
        .O(\rd_data[27]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[27]_i_14 
       (.I0(\rd_data[27]_i_28_n_0 ),
        .I1(\rd_data[27]_i_29_n_0 ),
        .I2(\rd_data[27]_i_30_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [27]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "rd_data[27]_i_14" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[27]_i_14_replica 
       (.I0(\rd_data[27]_i_28_n_0 ),
        .I1(\rd_data[27]_i_29_n_0 ),
        .I2(\rd_data[27]_i_30_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [27]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x[27]_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[27]_i_15 
       (.I0(\rd_data[27]_i_31_n_0 ),
        .I1(\rd_data[27]_i_32_n_0 ),
        .I2(\rd_data[27]_i_33_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [26]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[27]_i_16 
       (.I0(\rd_data[27]_i_34_n_0 ),
        .I1(\rd_data[27]_i_35_n_0 ),
        .I2(\rd_data[27]_i_36_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [25]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[27]_i_17 
       (.I0(\rd_data[27]_i_37_n_0 ),
        .I1(\rd_data[27]_i_38_n_0 ),
        .I2(\rd_data[27]_i_39_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [24]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[27]_i_18 
       (.I0(\processor/execute/alu_x [27]),
        .I1(\processor/execute/alu_y [27]),
        .O(\rd_data[27]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[27]_i_19 
       (.I0(\processor/execute/alu_x [26]),
        .I1(\processor/execute/alu_y [26]),
        .O(\rd_data[27]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[27]_i_2 
       (.I0(\rd_data[28]_i_4_n_0 ),
        .I1(\rd_data[27]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[27]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[28]_i_5_n_0 ),
        .O(\rd_data[27]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[27]_i_20 
       (.I0(\processor/execute/alu_x [25]),
        .I1(\processor/execute/alu_y [25]),
        .O(\rd_data[27]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[27]_i_21 
       (.I0(\processor/execute/alu_x [24]),
        .I1(\processor/execute/alu_y [24]),
        .O(\rd_data[27]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[27]_i_22 
       (.I0(\rd_data[27]_i_41_n_0 ),
        .I1(\csr_data_out[27]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [27]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \rd_data[27]_i_23 
       (.I0(\processor/execute/alu_x [31]),
        .I1(\processor/execute/alu_y [2]),
        .I2(\processor/execute/alu_y [4]),
        .I3(\processor/execute/alu_x [27]),
        .I4(\processor/execute/alu_y [3]),
        .O(\rd_data[27]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[27]_i_24 
       (.I0(\processor/execute/alu_x [27]),
        .I1(\processor/execute/alu_y [27]),
        .O(\rd_data[27]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[27]_i_25 
       (.I0(\processor/execute/alu_x [26]),
        .I1(\processor/execute/alu_y [26]),
        .O(\rd_data[27]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[27]_i_26 
       (.I0(\processor/execute/alu_x [25]),
        .I1(\processor/execute/alu_y [25]),
        .O(\rd_data[27]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[27]_i_27 
       (.I0(\processor/execute/alu_x [24]),
        .I1(\processor/execute/alu_y [24]),
        .O(\rd_data[27]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[27]_i_28 
       (.I0(\processor/ex_pc [27]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [27]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [27]),
        .O(\rd_data[27]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rd_data[27]_i_29 
       (.I0(\processor/mem_exception_context[badaddr] [27]),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .O(\rd_data[27]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[27]_i_3 
       (.I0(\rd_data[27]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [27]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[27]_i_8_n_0 ),
        .O(\rd_data[27]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000540455555555)) 
    \rd_data[27]_i_30 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\rd_data[27]_i_42_n_0 ),
        .I2(\csr_data_out[30]_i_9_n_0 ),
        .I3(\processor/wb_exception_context[badaddr] [27]),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\rd_data[27]_i_43_n_0 ),
        .O(\rd_data[27]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[27]_i_31 
       (.I0(\processor/ex_pc [26]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [26]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [26]),
        .O(\rd_data[27]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rd_data[27]_i_32 
       (.I0(\processor/mem_exception_context[badaddr] [26]),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .O(\rd_data[27]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000540455555555)) 
    \rd_data[27]_i_33 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\rd_data[27]_i_44_n_0 ),
        .I2(\csr_data_out[30]_i_9_n_0 ),
        .I3(\processor/wb_exception_context[badaddr] [26]),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\rd_data[27]_i_45_n_0 ),
        .O(\rd_data[27]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[27]_i_34 
       (.I0(\processor/ex_pc [25]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [25]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [25]),
        .O(\rd_data[27]_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rd_data[27]_i_35 
       (.I0(\processor/mem_exception_context[badaddr] [25]),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .O(\rd_data[27]_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000540455555555)) 
    \rd_data[27]_i_36 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\rd_data[27]_i_46_n_0 ),
        .I2(\csr_data_out[30]_i_9_n_0 ),
        .I3(\processor/wb_exception_context[badaddr] [25]),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\rd_data[27]_i_47_n_0 ),
        .O(\rd_data[27]_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[27]_i_37 
       (.I0(\processor/ex_pc [24]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [24]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [24]),
        .O(\rd_data[27]_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rd_data[27]_i_38 
       (.I0(\processor/mem_exception_context[badaddr] [24]),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .O(\rd_data[27]_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000540455555555)) 
    \rd_data[27]_i_39 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\rd_data[27]_i_48_n_0 ),
        .I2(\csr_data_out[30]_i_9_n_0 ),
        .I3(\processor/wb_exception_context[badaddr] [24]),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\rd_data[27]_i_49_n_0 ),
        .O(\rd_data[27]_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rd_data[27]_i_4 
       (.I0(\rd_data[27]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [1]),
        .I2(\rd_data[27]_i_10_n_0 ),
        .O(\rd_data[27]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[27]_i_41 
       (.I0(\processor/ex_pc [27]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [27]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [27]),
        .O(\rd_data[27]_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCAAACAAACAAAAAAA)) 
    \rd_data[27]_i_42 
       (.I0(\processor/csr_read_data [27]),
        .I1(\processor/wb_csr_data [27]),
        .I2(\processor/execute/csr_writeable ),
        .I3(\processor/execute/csr_value_forwarded3 ),
        .I4(\processor/wb_csr_write [1]),
        .I5(\processor/wb_csr_write [0]),
        .O(\rd_data[27]_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7F7F7FFF)) 
    \rd_data[27]_i_43 
       (.I0(\processor/mem_csr_data [27]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/mem_csr_write [0]),
        .I4(\processor/mem_csr_write [1]),
        .O(\rd_data[27]_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCAAACAAACAAAAAAA)) 
    \rd_data[27]_i_44 
       (.I0(\processor/csr_read_data [26]),
        .I1(\processor/wb_csr_data [26]),
        .I2(\processor/execute/csr_writeable ),
        .I3(\processor/execute/csr_value_forwarded3 ),
        .I4(\processor/wb_csr_write [1]),
        .I5(\processor/wb_csr_write [0]),
        .O(\rd_data[27]_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7F7F7FFF)) 
    \rd_data[27]_i_45 
       (.I0(\processor/mem_csr_data [26]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/mem_csr_write [0]),
        .I4(\processor/mem_csr_write [1]),
        .O(\rd_data[27]_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEAEAEAAA2A2A2AAA)) 
    \rd_data[27]_i_46 
       (.I0(\processor/csr_read_data [25]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded3 ),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/wb_csr_write [0]),
        .I5(\processor/wb_csr_data [25]),
        .O(\rd_data[27]_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7F7F7FFF)) 
    \rd_data[27]_i_47 
       (.I0(\processor/mem_csr_data [25]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/mem_csr_write [0]),
        .I4(\processor/mem_csr_write [1]),
        .O(\rd_data[27]_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEAEAEAAA2A2A2AAA)) 
    \rd_data[27]_i_48 
       (.I0(\processor/csr_read_data [24]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded3 ),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/wb_csr_write [0]),
        .I5(\processor/wb_csr_data [24]),
        .O(\rd_data[27]_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7F7F7FFF)) 
    \rd_data[27]_i_49 
       (.I0(\processor/mem_csr_data [24]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/mem_csr_write [0]),
        .I4(\processor/mem_csr_write [1]),
        .O(\rd_data[27]_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[27]_i_5 
       (.I0(\rd_data[29]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[31]_i_26_n_0 ),
        .I3(\rd_data[27]_i_11_n_0 ),
        .I4(\rd_data[31]_i_24_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[27]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[27]_i_6 
       (.I0(\rd_data[28]_i_11_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[27]_i_12_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [27]),
        .O(\rd_data[27]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[27]_i_8 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [27]),
        .I3(\processor/execute/alu_y [27]),
        .O(\rd_data[27]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF0F1F0E0)) 
    \rd_data[27]_i_9 
       (.I0(\processor/execute/alu_y [2]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [31]),
        .I3(\processor/execute/alu_y [4]),
        .I4(\processor/execute/alu_x [29]),
        .O(\rd_data[27]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[28]_i_1 
       (.I0(\rd_data[28]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[28]_i_3_n_0 ),
        .O(\processor/ex_rd_data [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h3300B8B8)) 
    \rd_data[28]_i_10 
       (.I0(\processor/execute/alu_x [5]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [21]),
        .I3(\processor/execute/alu_x [13]),
        .I4(\processor/execute/alu_y [3]),
        .O(\rd_data[28]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000B08)) 
    \rd_data[28]_i_11 
       (.I0(\processor/execute/alu_x [30]),
        .I1(\processor/execute/alu_y [1]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_x [28]),
        .I4(\processor/execute/alu_y [4]),
        .I5(\processor/execute/alu_y [2]),
        .O(\rd_data[28]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[28]_i_12 
       (.I0(\rd_data[28]_i_13_n_0 ),
        .I1(\csr_data_out[28]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [28]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[28]_i_13 
       (.I0(\processor/ex_pc [28]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [28]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [28]),
        .O(\rd_data[28]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[28]_i_2 
       (.I0(\rd_data[29]_i_4_n_0 ),
        .I1(\rd_data[28]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[28]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[29]_i_5_n_0 ),
        .O(\rd_data[28]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[28]_i_3 
       (.I0(\rd_data[28]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [28]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[28]_i_7_n_0 ),
        .O(\rd_data[28]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rd_data[28]_i_4 
       (.I0(\rd_data[28]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [1]),
        .I2(\rd_data[28]_i_9_n_0 ),
        .O(\rd_data[28]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[28]_i_5 
       (.I0(\rd_data[28]_i_10_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[31]_i_18_n_0 ),
        .I3(\rd_data[30]_i_12_n_0 ),
        .I4(\rd_data[31]_i_21_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[28]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[28]_i_6 
       (.I0(\rd_data[29]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[28]_i_11_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [28]),
        .O(\rd_data[28]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[28]_i_7 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [28]),
        .I3(\processor/execute/alu_y [28]),
        .O(\rd_data[28]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF0F1F0E0)) 
    \rd_data[28]_i_8 
       (.I0(\processor/execute/alu_y [2]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [31]),
        .I3(\processor/execute/alu_y [4]),
        .I4(\processor/execute/alu_x [30]),
        .O(\rd_data[28]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF0F1F0E0)) 
    \rd_data[28]_i_9 
       (.I0(\processor/execute/alu_y [2]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [31]),
        .I3(\processor/execute/alu_y [4]),
        .I4(\processor/execute/alu_x [28]),
        .O(\rd_data[28]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[29]_i_1 
       (.I0(\rd_data[29]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[29]_i_3_n_0 ),
        .O(\processor/ex_rd_data [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[29]_i_10 
       (.I0(\rd_data[29]_i_11_n_0 ),
        .I1(\csr_data_out[29]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [29]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[29]_i_11 
       (.I0(\processor/ex_pc [29]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [29]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [29]),
        .O(\rd_data[29]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[29]_i_2 
       (.I0(\rd_data[30]_i_4_n_0 ),
        .I1(\rd_data[29]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[29]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[30]_i_5_n_0 ),
        .O(\rd_data[29]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[29]_i_3 
       (.I0(\rd_data[29]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [29]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[29]_i_7_n_0 ),
        .O(\rd_data[29]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00FF01FF00FE00)) 
    \rd_data[29]_i_4 
       (.I0(\processor/execute/alu_y [1]),
        .I1(\processor/execute/alu_y [2]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_x [31]),
        .I4(\processor/execute/alu_y [4]),
        .I5(\processor/execute/alu_x [29]),
        .O(\rd_data[29]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[29]_i_5 
       (.I0(\rd_data[29]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[31]_i_26_n_0 ),
        .I3(\rd_data[31]_i_24_n_0 ),
        .I4(\rd_data[31]_i_25_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[29]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2F20FFFF2F200000)) 
    \rd_data[29]_i_6 
       (.I0(\rd_data[30]_i_13_n_0 ),
        .I1(\processor/execute/alu_y [1]),
        .I2(\processor/execute/alu_y [0]),
        .I3(\rd_data[29]_i_9_n_0 ),
        .I4(\processor/execute/alu_op [0]),
        .I5(\processor/execute/alu_instance/data6 [29]),
        .O(\rd_data[29]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[29]_i_7 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [29]),
        .I3(\processor/execute/alu_y [29]),
        .O(\rd_data[29]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h3300B8B8)) 
    \rd_data[29]_i_8 
       (.I0(\processor/execute/alu_x [6]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [22]),
        .I3(\processor/execute/alu_x [14]),
        .I4(\processor/execute/alu_y [3]),
        .O(\rd_data[29]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000B08)) 
    \rd_data[29]_i_9 
       (.I0(\processor/execute/alu_x [31]),
        .I1(\processor/execute/alu_y [1]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_x [29]),
        .I4(\processor/execute/alu_y [4]),
        .I5(\processor/execute/alu_y [2]),
        .O(\rd_data[29]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[2]_i_10 
       (.I0(\processor/ex_pc [2]),
        .I1(\processor/execute/shamt [2]),
        .I2(\processor/execute/alu_x_src [1]),
        .I3(\processor/execute/immediate [2]),
        .I4(\processor/execute/alu_x_src [0]),
        .I5(\processor/execute/rs1_forwarded [2]),
        .O(\rd_data[2]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[2]_i_12 
       (.I0(\processor/ex_pc [2]),
        .I1(\processor/execute/shamt [2]),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/immediate [2]),
        .I4(\processor/execute/alu_y_src [0]),
        .I5(\processor/ex_dmem_data_out [2]),
        .O(\rd_data[2]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rd_data[2]_i_14 
       (.I0(\rd_data[6]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[10]_i_12_n_0 ),
        .I3(\processor/execute/alu_y [3]),
        .I4(\rd_data[2]_i_23_n_0 ),
        .O(\rd_data[2]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rd_data[2]_i_17 
       (.I0(\processor/ex_pc [2]),
        .O(\rd_data[2]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8B8B8BB88BB88888)) 
    \rd_data[2]_i_2 
       (.I0(\rd_data[2]_i_4_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_x [2]),
        .I5(\processor/execute/alu_y [2]),
        .O(\rd_data[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rd_data[2]_i_21 
       (.I0(\processor/ex_pc [2]),
        .O(\rd_data[2]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rd_data[2]_i_23 
       (.I0(\processor/execute/alu_x [18]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [2]),
        .O(\rd_data[2]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \rd_data[2]_i_3 
       (.I0(\rd_data[3]_i_5_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[2]_i_7_n_0 ),
        .I3(\rd_data[31]_i_10_n_0 ),
        .I4(\processor/execute/alu_instance/data9 [2]),
        .I5(\rd_data[31]_i_11_n_0 ),
        .O(\rd_data[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \rd_data[2]_i_4 
       (.I0(\processor/execute/alu_instance/data7 [2]),
        .I1(\processor/execute/alu_instance/data6 [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data5 [2]),
        .O(\rd_data[2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[2]_i_5 
       (.I0(\rd_data[2]_i_10_n_0 ),
        .I1(\csr_data_out[2]_i_3_n_0 ),
        .I2(\processor/execute/alu_x_src [1]),
        .I3(\processor/execute/alu_x_src [2]),
        .I4(\processor/execute/alu_x_mux/data3 [2]),
        .I5(\processor/execute/alu_x_src [0]),
        .O(\processor/execute/alu_x [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h50CC50CC5FCC50CC)) 
    \rd_data[2]_i_6 
       (.I0(\csr_data_out[2]_i_3_n_0 ),
        .I1(\rd_data[2]_i_12_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [2]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \rd_data[2]_i_7 
       (.I0(\processor/execute/alu_y [2]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [1]),
        .I3(\processor/execute/alu_y [3]),
        .I4(\processor/execute/alu_y [1]),
        .O(\rd_data[2]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rd_data[2]_i_8 
       (.I0(\rd_data[3]_i_4_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[4]_i_8_n_0 ),
        .I3(\processor/execute/alu_y [1]),
        .I4(\rd_data[2]_i_14_n_0 ),
        .O(\processor/execute/alu_instance/data9 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rd_data[2]_i_9 
       (.I0(\rd_data[3]_i_11_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[4]_i_13_n_0 ),
        .I3(\processor/execute/alu_y [1]),
        .I4(\rd_data[2]_i_14_n_0 ),
        .O(\processor/execute/alu_instance/data7 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[30]_i_1 
       (.I0(\rd_data[30]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[30]_i_3_n_0 ),
        .O(\processor/ex_rd_data [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[30]_i_10 
       (.I0(\rd_data[30]_i_25_n_0 ),
        .I1(\csr_data_out[4]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [4]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[30]_i_11 
       (.I0(\rd_data[30]_i_26_n_0 ),
        .I1(\rd_data[30]_i_27_n_0 ),
        .I2(\rd_data[30]_i_28_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [30]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h3300B8B8)) 
    \rd_data[30]_i_12 
       (.I0(\processor/execute/alu_x [7]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [23]),
        .I3(\processor/execute/alu_x [15]),
        .I4(\processor/execute/alu_y [3]),
        .O(\rd_data[30]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \rd_data[30]_i_13 
       (.I0(\processor/execute/alu_y [3]),
        .I1(\processor/execute/alu_x [30]),
        .I2(\processor/execute/alu_y [4]),
        .I3(\processor/execute/alu_y [2]),
        .O(\rd_data[30]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[30]_i_14 
       (.I0(\rd_data[30]_i_31_n_0 ),
        .I1(\rd_data[30]_i_32_n_0 ),
        .I2(\rd_data[30]_i_33_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [29]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[30]_i_15 
       (.I0(\rd_data[30]_i_34_n_0 ),
        .I1(\rd_data[30]_i_35_n_0 ),
        .I2(\rd_data[30]_i_36_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [28]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[30]_i_16 
       (.I0(\processor/execute/alu_y [31]),
        .I1(\processor/execute/alu_x [31]),
        .O(\rd_data[30]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[30]_i_17 
       (.I0(\processor/execute/alu_x [30]),
        .I1(\processor/execute/alu_y [30]),
        .O(\rd_data[30]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[30]_i_18 
       (.I0(\processor/execute/alu_x [29]),
        .I1(\processor/execute/alu_y [29]),
        .O(\rd_data[30]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[30]_i_19 
       (.I0(\processor/execute/alu_x [28]),
        .I1(\processor/execute/alu_y [28]),
        .O(\rd_data[30]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[30]_i_2 
       (.I0(\processor/execute/alu_x [31]),
        .I1(\rd_data[30]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[30]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[31]_i_9_n_0 ),
        .O(\rd_data[30]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[30]_i_20 
       (.I0(\rd_data[30]_i_37_n_0 ),
        .I1(\csr_data_out[30]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [30]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[30]_i_21 
       (.I0(\processor/ex_pc [3]),
        .I1(\processor/execute/shamt [3]),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/immediate [3]),
        .I4(\processor/execute/alu_y_src [0]),
        .I5(\processor/ex_dmem_data_out [3]),
        .O(\rd_data[30]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000EFEF00EF)) 
    \rd_data[30]_i_22 
       (.I0(\rd_data[30]_i_38_n_0 ),
        .I1(\csr_data_out[3]_i_8_n_0 ),
        .I2(\rd_data[30]_i_39_n_0 ),
        .I3(\rd_data[30]_i_40_n_0 ),
        .I4(\rd_data[30]_i_41_n_0 ),
        .I5(\csr_data_out[31]_i_6_n_0 ),
        .O(\rd_data[30]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \rd_data[30]_i_23 
       (.I0(\processor/execute/alu_y_src [1]),
        .I1(\processor/execute/alu_y_src [2]),
        .O(\rd_data[30]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h5D)) 
    \rd_data[30]_i_24 
       (.I0(\processor/execute/alu_y_src [2]),
        .I1(\processor/execute/alu_y_src [0]),
        .I2(\processor/execute/alu_y_src [1]),
        .O(\rd_data[30]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[30]_i_25 
       (.I0(\processor/ex_pc [4]),
        .I1(\processor/execute/shamt [4]),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/immediate [4]),
        .I4(\processor/execute/alu_y_src [0]),
        .I5(\processor/ex_dmem_data_out [4]),
        .O(\rd_data[30]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[30]_i_26 
       (.I0(\processor/ex_pc [30]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [30]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [30]),
        .O(\rd_data[30]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rd_data[30]_i_27 
       (.I0(\processor/mem_exception_context[badaddr] [30]),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .O(\rd_data[30]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000540455555555)) 
    \rd_data[30]_i_28 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\rd_data[30]_i_42_n_0 ),
        .I2(\csr_data_out[30]_i_9_n_0 ),
        .I3(\processor/wb_exception_context[badaddr] [30]),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\rd_data[30]_i_43_n_0 ),
        .O(\rd_data[30]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \rd_data[30]_i_29 
       (.I0(\processor/execute/alu_x_src [1]),
        .I1(\processor/execute/alu_x_src [2]),
        .O(\rd_data[30]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[30]_i_3 
       (.I0(\rd_data[30]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [30]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[30]_i_8_n_0 ),
        .O(\rd_data[30]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h5D)) 
    \rd_data[30]_i_30 
       (.I0(\processor/execute/alu_x_src [2]),
        .I1(\processor/execute/alu_x_src [0]),
        .I2(\processor/execute/alu_x_src [1]),
        .O(\rd_data[30]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[30]_i_31 
       (.I0(\processor/ex_pc [29]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [29]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [29]),
        .O(\rd_data[30]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rd_data[30]_i_32 
       (.I0(\processor/mem_exception_context[badaddr] [29]),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .O(\rd_data[30]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000540455555555)) 
    \rd_data[30]_i_33 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\rd_data[30]_i_44_n_0 ),
        .I2(\csr_data_out[30]_i_9_n_0 ),
        .I3(\processor/wb_exception_context[badaddr] [29]),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\rd_data[30]_i_45_n_0 ),
        .O(\rd_data[30]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[30]_i_34 
       (.I0(\processor/ex_pc [28]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [28]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [28]),
        .O(\rd_data[30]_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rd_data[30]_i_35 
       (.I0(\processor/mem_exception_context[badaddr] [28]),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .O(\rd_data[30]_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000540455555555)) 
    \rd_data[30]_i_36 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\rd_data[30]_i_46_n_0 ),
        .I2(\csr_data_out[30]_i_9_n_0 ),
        .I3(\processor/wb_exception_context[badaddr] [28]),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\rd_data[30]_i_47_n_0 ),
        .O(\rd_data[30]_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[30]_i_37 
       (.I0(\processor/ex_pc [30]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [30]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [30]),
        .O(\rd_data[30]_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2000202020202020)) 
    \rd_data[30]_i_38 
       (.I0(\processor/wb_exception_context ),
        .I1(\rd_data[30]_i_48_n_0 ),
        .I2(\processor/wb_exception ),
        .I3(\csr_data_out[31]_i_18_n_0 ),
        .I4(\processor/execute/csr_value_forwarded30_out ),
        .I5(\processor/execute/csr_writeable ),
        .O(\rd_data[30]_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD0DDDDDDDFDDDDDD)) 
    \rd_data[30]_i_39 
       (.I0(\csr_data_out[31]_i_16_n_0 ),
        .I1(\csr_data_out[31]_i_19_n_0 ),
        .I2(\csr_data_out[31]_i_18_n_0 ),
        .I3(\processor/execute/csr_value_forwarded30_out ),
        .I4(\processor/execute/csr_writeable ),
        .I5(\processor/mem_csr_data [3]),
        .O(\rd_data[30]_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00FF01FF00FE00)) 
    \rd_data[30]_i_4 
       (.I0(\processor/execute/alu_y [1]),
        .I1(\processor/execute/alu_y [2]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_x [31]),
        .I4(\processor/execute/alu_y [4]),
        .I5(\processor/execute/alu_x [30]),
        .O(\rd_data[30]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h57777777F7777777)) 
    \rd_data[30]_i_40 
       (.I0(\csr_data_out[31]_i_21_n_0 ),
        .I1(\processor/csr_read_data [3]),
        .I2(\processor/csr_unit/tohost_data1__0 ),
        .I3(\processor/execute/csr_value_forwarded3 ),
        .I4(\processor/execute/csr_writeable ),
        .I5(\processor/wb_csr_data [3]),
        .O(\rd_data[30]_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF55D5)) 
    \rd_data[30]_i_41 
       (.I0(\csr_data_out[31]_i_16_n_0 ),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\csr_data_out[31]_i_18_n_0 ),
        .I4(\csr_data_out[31]_i_19_n_0 ),
        .I5(\rd_data[30]_i_49_n_0 ),
        .O(\rd_data[30]_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCAAACAAACAAAAAAA)) 
    \rd_data[30]_i_42 
       (.I0(\processor/csr_read_data [30]),
        .I1(\processor/wb_csr_data [30]),
        .I2(\processor/execute/csr_writeable ),
        .I3(\processor/execute/csr_value_forwarded3 ),
        .I4(\processor/wb_csr_write [1]),
        .I5(\processor/wb_csr_write [0]),
        .O(\rd_data[30]_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7F7F7FFF)) 
    \rd_data[30]_i_43 
       (.I0(\processor/mem_csr_data [30]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/mem_csr_write [0]),
        .I4(\processor/mem_csr_write [1]),
        .O(\rd_data[30]_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEAEAEAAA2A2A2AAA)) 
    \rd_data[30]_i_44 
       (.I0(\processor/csr_read_data [29]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded3 ),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/wb_csr_write [0]),
        .I5(\processor/wb_csr_data [29]),
        .O(\rd_data[30]_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7F7F7FFF)) 
    \rd_data[30]_i_45 
       (.I0(\processor/mem_csr_data [29]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/mem_csr_write [0]),
        .I4(\processor/mem_csr_write [1]),
        .O(\rd_data[30]_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCAAACAAACAAAAAAA)) 
    \rd_data[30]_i_46 
       (.I0(\processor/csr_read_data [28]),
        .I1(\processor/wb_csr_data [28]),
        .I2(\processor/execute/csr_writeable ),
        .I3(\processor/execute/csr_value_forwarded3 ),
        .I4(\processor/wb_csr_write [1]),
        .I5(\processor/wb_csr_write [0]),
        .O(\rd_data[30]_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7F7F7FFF)) 
    \rd_data[30]_i_47 
       (.I0(\processor/mem_csr_data [28]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/mem_csr_write [0]),
        .I4(\processor/mem_csr_write [1]),
        .O(\rd_data[30]_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rd_data[30]_i_48 
       (.I0(\csr_data_out[11]_i_8_n_0 ),
        .I1(\rd_data[30]_i_50_n_0 ),
        .I2(\processor/ex_csr_address [4]),
        .I3(\csr_data_out[30]_i_11_n_0 ),
        .I4(\processor/ex_csr_address [5]),
        .I5(\processor/ex_csr_address[3]_repN ),
        .O(\rd_data[30]_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \rd_data[30]_i_49 
       (.I0(\processor/wb_exception_context[badaddr] [3]),
        .I1(\processor/wb_exception ),
        .I2(\csr_data_out[31]_i_14_n_0 ),
        .I3(\csr_data_out[31]_i_15_n_0 ),
        .I4(\csr_data_out[31]_i_31_n_0 ),
        .I5(\processor/ex_csr_address [0]),
        .O(\rd_data[30]_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[30]_i_5 
       (.I0(\rd_data[30]_i_12_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[31]_i_21_n_0 ),
        .I3(\rd_data[31]_i_18_n_0 ),
        .I4(\rd_data[31]_i_19_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[30]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \rd_data[30]_i_50 
       (.I0(\processor/ex_csr_address [9]),
        .I1(\processor/ex_csr_address [8]),
        .O(\rd_data[30]_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF022FFFFF0220000)) 
    \rd_data[30]_i_6 
       (.I0(\rd_data[30]_i_13_n_0 ),
        .I1(\processor/execute/alu_y [1]),
        .I2(\rd_data[31]_i_12_n_0 ),
        .I3(\processor/execute/alu_y [0]),
        .I4(\processor/execute/alu_op [0]),
        .I5(\processor/execute/alu_instance/data6 [30]),
        .O(\rd_data[30]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[30]_i_8 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [30]),
        .I3(\processor/execute/alu_y [30]),
        .O(\rd_data[30]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[30]_i_9 
       (.I0(\rd_data[30]_i_21_n_0 ),
        .I1(\csr_data_out[3]_i_7_n_0 ),
        .I2(\rd_data[30]_i_22_n_0 ),
        .I3(\rd_data[30]_i_23_n_0 ),
        .I4(\processor/execute/alu_y_mux/data3 [3]),
        .I5(\rd_data[30]_i_24_n_0 ),
        .O(\processor/execute/alu_y [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBA)) 
    \rd_data[31]_i_10 
       (.I0(\processor/execute/alu_op [2]),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .O(\rd_data[31]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \rd_data[31]_i_11 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [2]),
        .O(\rd_data[31]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \rd_data[31]_i_12 
       (.I0(\processor/execute/alu_y [2]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [31]),
        .I3(\processor/execute/alu_y [3]),
        .I4(\processor/execute/alu_y [1]),
        .O(\rd_data[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[31]_i_14 
       (.I0(\processor/ex_pc [31]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [31]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [31]),
        .O(\rd_data[31]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[31]_i_16 
       (.I0(\processor/ex_pc [31]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [31]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [31]),
        .O(\rd_data[31]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \rd_data[31]_i_18 
       (.I0(\processor/execute/alu_x [1]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [17]),
        .I3(\processor/execute/alu_y [3]),
        .I4(\processor/execute/alu_x [9]),
        .I5(\processor/execute/alu_x [25]),
        .O(\rd_data[31]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \rd_data[31]_i_19 
       (.I0(\processor/execute/alu_x [5]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [21]),
        .I3(\processor/execute/alu_y [3]),
        .I4(\processor/execute/alu_x [13]),
        .I5(\processor/execute/alu_x [29]),
        .O(\rd_data[31]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8B8B8BB88BB88888)) 
    \rd_data[31]_i_2 
       (.I0(\rd_data[31]_i_4_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_x [31]),
        .I5(\processor/execute/alu_y [31]),
        .O(\rd_data[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h50CC50CC5FCC50CC)) 
    \rd_data[31]_i_20 
       (.I0(\csr_data_out[1]_i_3_n_0 ),
        .I1(\rd_data[31]_i_40_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [1]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \rd_data[31]_i_21 
       (.I0(\processor/execute/alu_x [3]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [19]),
        .I3(\processor/execute/alu_y [3]),
        .I4(\processor/execute/alu_x [11]),
        .I5(\processor/execute/alu_x [27]),
        .O(\rd_data[31]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \rd_data[31]_i_22 
       (.I0(\processor/execute/alu_x [7]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [23]),
        .I3(\processor/execute/alu_y [3]),
        .I4(\processor/execute/alu_x [15]),
        .I5(\processor/execute/alu_x [31]),
        .O(\rd_data[31]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[31]_i_23 
       (.I0(\processor/ex_pc [0]),
        .I1(\processor/execute/shamt [0]),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/immediate [0]),
        .I4(\processor/execute/alu_y_src [0]),
        .I5(\processor/ex_dmem_data_out [0]),
        .O(\rd_data[31]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \rd_data[31]_i_24 
       (.I0(\processor/execute/alu_x [0]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [16]),
        .I3(\processor/execute/alu_y [3]),
        .I4(\processor/execute/alu_x [8]),
        .I5(\processor/execute/alu_x [24]),
        .O(\rd_data[31]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \rd_data[31]_i_25 
       (.I0(\processor/execute/alu_x [4]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [20]),
        .I3(\processor/execute/alu_y [3]),
        .I4(\processor/execute/alu_x [12]),
        .I5(\processor/execute/alu_x [28]),
        .O(\rd_data[31]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \rd_data[31]_i_26 
       (.I0(\processor/execute/alu_x [2]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [18]),
        .I3(\processor/execute/alu_y [3]),
        .I4(\processor/execute/alu_x [10]),
        .I5(\processor/execute/alu_x [26]),
        .O(\rd_data[31]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \rd_data[31]_i_27 
       (.I0(\processor/execute/alu_x [6]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [22]),
        .I3(\processor/execute/alu_y [3]),
        .I4(\processor/execute/alu_x [14]),
        .I5(\processor/execute/alu_x [30]),
        .O(\rd_data[31]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[31]_i_28 
       (.I0(\processor/execute/alu_x [31]),
        .I1(\processor/execute/alu_y [31]),
        .O(\rd_data[31]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[31]_i_29 
       (.I0(\processor/execute/alu_x [30]),
        .I1(\processor/execute/alu_y [30]),
        .O(\rd_data[31]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \rd_data[31]_i_3 
       (.I0(\rd_data[31]_i_7_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[31]_i_9_n_0 ),
        .I3(\rd_data[31]_i_10_n_0 ),
        .I4(\processor/execute/alu_x [31]),
        .I5(\rd_data[31]_i_11_n_0 ),
        .O(\rd_data[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[31]_i_30 
       (.I0(\processor/execute/alu_x [29]),
        .I1(\processor/execute/alu_y [29]),
        .O(\rd_data[31]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[31]_i_31 
       (.I0(\processor/execute/alu_x [28]),
        .I1(\processor/execute/alu_y [28]),
        .O(\rd_data[31]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h22FFF0002200F000)) 
    \rd_data[31]_i_4 
       (.I0(\rd_data[31]_i_12_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\processor/execute/alu_instance/data6 [31]),
        .I3(\processor/execute/alu_op [1]),
        .I4(\processor/execute/alu_op [0]),
        .I5(\processor/execute/alu_instance/data5 [31]),
        .O(\rd_data[31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[31]_i_40 
       (.I0(\processor/ex_pc [1]),
        .I1(\processor/execute/shamt [1]),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/immediate [1]),
        .I4(\processor/execute/alu_y_src [0]),
        .I5(\processor/ex_dmem_data_out [1]),
        .O(\rd_data[31]_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[31]_i_5 
       (.I0(\rd_data[31]_i_14_n_0 ),
        .I1(\csr_data_out[31]_i_4_n_0 ),
        .I2(\processor/execute/alu_x_src [1]),
        .I3(\processor/execute/alu_x_src [2]),
        .I4(\processor/execute/alu_x_mux/data3 [31]),
        .I5(\processor/execute/alu_x_src [0]),
        .O(\processor/execute/alu_x [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h50CC50CC5FCC50CC)) 
    \rd_data[31]_i_6 
       (.I0(\csr_data_out[31]_i_4_n_0 ),
        .I1(\rd_data[31]_i_16_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [31]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \rd_data[31]_i_7 
       (.I0(\rd_data[31]_i_18_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[31]_i_19_n_0 ),
        .I3(\processor/execute/alu_y [1]),
        .I4(\rd_data[31]_i_21_n_0 ),
        .I5(\rd_data[31]_i_22_n_0 ),
        .O(\rd_data[31]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[31]_i_8 
       (.I0(\rd_data[31]_i_23_n_0 ),
        .I1(\csr_data_out[0]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/ex_pc [0]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \rd_data[31]_i_9 
       (.I0(\rd_data[31]_i_24_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[31]_i_25_n_0 ),
        .I3(\processor/execute/alu_y [1]),
        .I4(\rd_data[31]_i_26_n_0 ),
        .I5(\rd_data[31]_i_27_n_0 ),
        .O(\rd_data[31]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[3]_i_1 
       (.I0(\rd_data[3]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[3]_i_3_n_0 ),
        .O(\processor/ex_rd_data [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00CFFFCF00)) 
    \rd_data[3]_i_10 
       (.I0(\rd_data[3]_i_19_n_0 ),
        .I1(\csr_data_out[0]_i_7_n_0 ),
        .I2(\rd_data[3]_i_20_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/ex_pc [0]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[3]_i_11 
       (.I0(\rd_data[9]_i_12_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[5]_i_8_n_0 ),
        .I3(\processor/execute/alu_y [1]),
        .I4(\rd_data[3]_i_9_n_0 ),
        .O(\rd_data[3]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[3]_i_13 
       (.I0(\rd_data[3]_i_25_n_0 ),
        .I1(\csr_data_out[3]_i_7_n_0 ),
        .I2(\rd_data[30]_i_22_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [3]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[3]_i_14 
       (.I0(\processor/execute/alu_x [3]),
        .I1(\processor/execute/alu_y [3]),
        .O(\rd_data[3]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[3]_i_15 
       (.I0(\processor/execute/alu_x [2]),
        .I1(\processor/execute/alu_y [2]),
        .O(\rd_data[3]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[3]_i_16 
       (.I0(\processor/execute/alu_x [1]),
        .I1(\processor/execute/alu_y [1]),
        .O(\rd_data[3]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[3]_i_17 
       (.I0(\processor/execute/alu_x [0]),
        .I1(\processor/execute/alu_y [0]),
        .O(\rd_data[3]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rd_data[3]_i_18 
       (.I0(\processor/execute/alu_x [19]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [3]),
        .O(\rd_data[3]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[3]_i_19 
       (.I0(\processor/ex_pc [0]),
        .I1(\processor/execute/shamt [0]),
        .I2(\processor/execute/alu_x_src [1]),
        .I3(\processor/execute/immediate [0]),
        .I4(\processor/execute/alu_x_src [0]),
        .I5(\processor/execute/rs1_forwarded [0]),
        .O(\rd_data[3]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[3]_i_2 
       (.I0(\rd_data[4]_i_4_n_0 ),
        .I1(\rd_data[3]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[3]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[4]_i_5_n_0 ),
        .O(\rd_data[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF444400F0)) 
    \rd_data[3]_i_20 
       (.I0(\rd_data[3]_i_26_n_0 ),
        .I1(\rd_data[3]_i_27_n_0 ),
        .I2(\rd_data[3]_i_28_n_0 ),
        .I3(\rd_data[3]_i_29_n_0 ),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\csr_data_out[31]_i_6_n_0 ),
        .O(\rd_data[3]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[3]_i_21 
       (.I0(\processor/execute/alu_x [3]),
        .I1(\processor/execute/alu_y [3]),
        .O(\rd_data[3]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[3]_i_22 
       (.I0(\processor/execute/alu_x [2]),
        .I1(\processor/execute/alu_y [2]),
        .O(\rd_data[3]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[3]_i_23 
       (.I0(\processor/execute/alu_x [1]),
        .I1(\processor/execute/alu_y [1]),
        .O(\rd_data[3]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[3]_i_24 
       (.I0(\processor/execute/alu_x [0]),
        .I1(\processor/execute/alu_y [0]),
        .O(\rd_data[3]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[3]_i_25 
       (.I0(\processor/ex_pc [3]),
        .I1(\processor/execute/shamt [3]),
        .I2(\processor/execute/alu_x_src [1]),
        .I3(\processor/execute/immediate [3]),
        .I4(\processor/execute/alu_x_src [0]),
        .I5(\processor/execute/rs1_forwarded [3]),
        .O(\rd_data[3]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2000202020202020)) 
    \rd_data[3]_i_26 
       (.I0(\processor/wb_exception_context[ie] ),
        .I1(\rd_data[30]_i_48_n_0 ),
        .I2(\processor/wb_exception ),
        .I3(\csr_data_out[31]_i_18_n_0 ),
        .I4(\processor/execute/csr_value_forwarded30_out ),
        .I5(\processor/execute/csr_writeable ),
        .O(\rd_data[3]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCF55CFCFCFCFCFCF)) 
    \rd_data[3]_i_27 
       (.I0(\processor/mem_csr_data [0]),
        .I1(\csr_data_out[3]_i_10_n_0 ),
        .I2(\processor/wb_exception_context[cause] [0]),
        .I3(\csr_data_out[31]_i_18_n_0 ),
        .I4(\processor/execute/csr_value_forwarded30_out ),
        .I5(\processor/execute/csr_writeable ),
        .O(\rd_data[3]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h57777777F7777777)) 
    \rd_data[3]_i_28 
       (.I0(\csr_data_out[31]_i_21_n_0 ),
        .I1(\processor/csr_read_data [0]),
        .I2(\processor/csr_unit/tohost_data1__0 ),
        .I3(\processor/execute/csr_value_forwarded3 ),
        .I4(\processor/execute/csr_writeable ),
        .I5(\processor/wb_csr_data [0]),
        .O(\rd_data[3]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \rd_data[3]_i_29 
       (.I0(\processor/wb_exception_context[badaddr] [0]),
        .I1(\csr_data_out[31]_i_21_n_0 ),
        .O(\rd_data[3]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[3]_i_3 
       (.I0(\rd_data[3]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [3]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[3]_i_8_n_0 ),
        .O(\rd_data[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[3]_i_4 
       (.I0(\rd_data[9]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[5]_i_8_n_0 ),
        .I3(\processor/execute/alu_y [1]),
        .I4(\rd_data[3]_i_9_n_0 ),
        .O(\rd_data[3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000002030200)) 
    \rd_data[3]_i_5 
       (.I0(\processor/execute/alu_x [0]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_y [1]),
        .I4(\processor/execute/alu_x [2]),
        .I5(\processor/execute/alu_y [2]),
        .O(\rd_data[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[3]_i_6 
       (.I0(\rd_data[4]_i_10_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[3]_i_11_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [3]),
        .O(\rd_data[3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[3]_i_8 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [3]),
        .I3(\processor/execute/alu_y [3]),
        .O(\rd_data[3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rd_data[3]_i_9 
       (.I0(\rd_data[7]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[11]_i_22_n_0 ),
        .I3(\processor/execute/alu_y [3]),
        .I4(\rd_data[3]_i_18_n_0 ),
        .O(\rd_data[3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[4]_i_1 
       (.I0(\rd_data[4]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[4]_i_3_n_0 ),
        .O(\processor/ex_rd_data [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[4]_i_10 
       (.I0(\rd_data[10]_i_13_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[6]_i_8_n_0 ),
        .I3(\processor/execute/alu_y [1]),
        .I4(\rd_data[4]_i_13_n_0 ),
        .O(\rd_data[4]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[4]_i_11 
       (.I0(\processor/execute/alu_x [28]),
        .I1(\processor/execute/alu_x [12]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_x [20]),
        .I4(\processor/execute/alu_y [4]),
        .I5(\processor/execute/alu_x [4]),
        .O(\rd_data[4]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[4]_i_12 
       (.I0(\processor/ex_pc [1]),
        .I1(\processor/execute/shamt [1]),
        .I2(\processor/execute/alu_x_src [1]),
        .I3(\processor/execute/immediate [1]),
        .I4(\processor/execute/alu_x_src [0]),
        .I5(\processor/execute/rs1_forwarded [1]),
        .O(\rd_data[4]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rd_data[4]_i_13 
       (.I0(\rd_data[8]_i_12_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[4]_i_11_n_0 ),
        .O(\rd_data[4]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[4]_i_2 
       (.I0(\rd_data[5]_i_4_n_0 ),
        .I1(\rd_data[4]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[4]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[5]_i_5_n_0 ),
        .O(\rd_data[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[4]_i_3 
       (.I0(\rd_data[4]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [4]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[4]_i_7_n_0 ),
        .O(\rd_data[4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[4]_i_4 
       (.I0(\rd_data[10]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[6]_i_8_n_0 ),
        .I3(\processor/execute/alu_y [1]),
        .I4(\rd_data[4]_i_8_n_0 ),
        .O(\rd_data[4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000030022222222)) 
    \rd_data[4]_i_5 
       (.I0(\rd_data[10]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_x [1]),
        .I4(\processor/execute/alu_y [4]),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[4]_i_6 
       (.I0(\rd_data[5]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[4]_i_10_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [4]),
        .O(\rd_data[4]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[4]_i_7 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [4]),
        .I3(\processor/execute/alu_y [4]),
        .O(\rd_data[4]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rd_data[4]_i_8 
       (.I0(\rd_data[8]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[4]_i_11_n_0 ),
        .O(\rd_data[4]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "rd_data[4]_i_8" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rd_data[4]_i_8_replica 
       (.I0(\rd_data[8]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[4]_i_11_n_0 ),
        .O(\rd_data[4]_i_8_n_0_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[4]_i_9 
       (.I0(\rd_data[4]_i_12_n_0 ),
        .I1(\csr_data_out[1]_i_3_n_0 ),
        .I2(\processor/execute/alu_x_src [1]),
        .I3(\processor/execute/alu_x_src [2]),
        .I4(\processor/execute/alu_x_mux/data3 [1]),
        .I5(\processor/execute/alu_x_src [0]),
        .O(\processor/execute/alu_x [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[5]_i_1 
       (.I0(\rd_data[5]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[5]_i_3_n_0 ),
        .O(\processor/ex_rd_data [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[5]_i_10 
       (.I0(\rd_data[5]_i_11_n_0 ),
        .I1(\csr_data_out[5]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [5]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[5]_i_11 
       (.I0(\processor/ex_pc [5]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [5]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [5]),
        .O(\rd_data[5]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[5]_i_2 
       (.I0(\rd_data[6]_i_4_n_0 ),
        .I1(\rd_data[5]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[5]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[6]_i_5_n_0 ),
        .O(\rd_data[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[5]_i_3 
       (.I0(\rd_data[5]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [5]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[5]_i_7_n_0 ),
        .O(\rd_data[5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[5]_i_4 
       (.I0(\rd_data[9]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[5]_i_8_n_0 ),
        .I3(\rd_data[11]_i_9_n_0 ),
        .I4(\rd_data[7]_i_9_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[5]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \rd_data[5]_i_5 
       (.I0(\processor/execute/alu_y [3]),
        .I1(\processor/execute/alu_x [2]),
        .I2(\processor/execute/alu_y [4]),
        .I3(\processor/execute/alu_y [2]),
        .I4(\processor/execute/alu_y [1]),
        .I5(\rd_data[7]_i_10_n_0 ),
        .O(\rd_data[5]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[5]_i_6 
       (.I0(\rd_data[6]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[5]_i_9_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [5]),
        .O(\rd_data[5]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[5]_i_7 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [5]),
        .I3(\processor/execute/alu_y [5]),
        .O(\rd_data[5]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[5]_i_8 
       (.I0(\processor/execute/alu_x [29]),
        .I1(\processor/execute/alu_x [13]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_x [21]),
        .I4(\processor/execute/alu_y [4]),
        .I5(\processor/execute/alu_x [5]),
        .O(\rd_data[5]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[5]_i_9 
       (.I0(\rd_data[9]_i_12_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[5]_i_8_n_0 ),
        .I3(\rd_data[11]_i_23_n_0 ),
        .I4(\rd_data[7]_i_9_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[5]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[6]_i_1 
       (.I0(\rd_data[6]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[6]_i_3_n_0 ),
        .O(\processor/ex_rd_data [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[6]_i_10 
       (.I0(\rd_data[6]_i_11_n_0 ),
        .I1(\csr_data_out[6]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [6]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[6]_i_11 
       (.I0(\processor/ex_pc [6]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [6]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [6]),
        .O(\rd_data[6]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[6]_i_2 
       (.I0(\rd_data[7]_i_4_n_0 ),
        .I1(\rd_data[6]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[6]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[7]_i_5_n_0 ),
        .O(\rd_data[6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[6]_i_3 
       (.I0(\rd_data[6]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [6]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[6]_i_7_n_0 ),
        .O(\rd_data[6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[6]_i_4 
       (.I0(\rd_data[10]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[6]_i_8_n_0 ),
        .I3(\rd_data[12]_i_8_n_0 ),
        .I4(\rd_data[8]_i_8_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[6]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \rd_data[6]_i_5 
       (.I0(\rd_data[10]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\processor/execute/alu_y [1]),
        .I3(\rd_data[8]_i_9_n_0 ),
        .O(\rd_data[6]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[6]_i_6 
       (.I0(\rd_data[7]_i_11_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[6]_i_9_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [6]),
        .O(\rd_data[6]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[6]_i_7 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [6]),
        .I3(\processor/execute/alu_y [6]),
        .O(\rd_data[6]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[6]_i_8 
       (.I0(\processor/execute/alu_x [30]),
        .I1(\processor/execute/alu_x [14]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_x [22]),
        .I4(\processor/execute/alu_y [4]),
        .I5(\processor/execute/alu_x [6]),
        .O(\rd_data[6]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[6]_i_9 
       (.I0(\rd_data[12]_i_12_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[8]_i_12_n_0 ),
        .I3(\rd_data[10]_i_13_n_0 ),
        .I4(\rd_data[6]_i_8_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[6]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[7]_i_1 
       (.I0(\rd_data[7]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[7]_i_3_n_0 ),
        .O(\processor/ex_rd_data [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02030200)) 
    \rd_data[7]_i_10 
       (.I0(\processor/execute/alu_x [0]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_y [2]),
        .I4(\processor/execute/alu_x [4]),
        .O(\rd_data[7]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[7]_i_11 
       (.I0(\rd_data[13]_i_12_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[9]_i_12_n_0 ),
        .I3(\rd_data[11]_i_23_n_0 ),
        .I4(\rd_data[7]_i_9_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[7]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[7]_i_13 
       (.I0(\rd_data[7]_i_26_n_0 ),
        .I1(\rd_data[7]_i_27_n_0 ),
        .I2(\rd_data[7]_i_28_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [7]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[7]_i_14 
       (.I0(\rd_data[7]_i_29_n_0 ),
        .I1(\rd_data[7]_i_30_n_0 ),
        .I2(\rd_data[7]_i_31_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [6]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00FCFFFC00)) 
    \rd_data[7]_i_15 
       (.I0(\rd_data[7]_i_32_n_0 ),
        .I1(\rd_data[7]_i_33_n_0 ),
        .I2(\rd_data[7]_i_34_n_0 ),
        .I3(\rd_data[30]_i_29_n_0 ),
        .I4(\processor/execute/alu_x_mux/data3 [5]),
        .I5(\rd_data[30]_i_30_n_0 ),
        .O(\processor/execute/alu_x [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[7]_i_16 
       (.I0(\rd_data[7]_i_35_n_0 ),
        .I1(\csr_data_out[4]_i_3_n_0 ),
        .I2(\processor/execute/alu_x_src [1]),
        .I3(\processor/execute/alu_x_src [2]),
        .I4(\processor/execute/alu_x_mux/data3 [4]),
        .I5(\processor/execute/alu_x_src [0]),
        .O(\processor/execute/alu_x [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[7]_i_17 
       (.I0(\processor/execute/alu_x [7]),
        .I1(\processor/execute/alu_y [7]),
        .O(\rd_data[7]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[7]_i_18 
       (.I0(\processor/execute/alu_x [6]),
        .I1(\processor/execute/alu_y [6]),
        .O(\rd_data[7]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[7]_i_19 
       (.I0(\processor/execute/alu_x [5]),
        .I1(\processor/execute/alu_y [5]),
        .O(\rd_data[7]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[7]_i_2 
       (.I0(\rd_data[8]_i_4_n_0 ),
        .I1(\rd_data[7]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[7]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[8]_i_5_n_0 ),
        .O(\rd_data[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rd_data[7]_i_20 
       (.I0(\processor/execute/alu_x [4]),
        .I1(\processor/execute/alu_y [4]),
        .O(\rd_data[7]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[7]_i_21 
       (.I0(\rd_data[7]_i_36_n_0 ),
        .I1(\csr_data_out[7]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [7]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[7]_i_22 
       (.I0(\processor/execute/alu_x [7]),
        .I1(\processor/execute/alu_y [7]),
        .O(\rd_data[7]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[7]_i_23 
       (.I0(\processor/execute/alu_x [6]),
        .I1(\processor/execute/alu_y [6]),
        .O(\rd_data[7]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[7]_i_24 
       (.I0(\processor/execute/alu_x [5]),
        .I1(\processor/execute/alu_y [5]),
        .O(\rd_data[7]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \rd_data[7]_i_25 
       (.I0(\processor/execute/alu_x [4]),
        .I1(\processor/execute/alu_y [4]),
        .O(\rd_data[7]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[7]_i_26 
       (.I0(\processor/ex_pc [7]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [7]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded[7]_repN ),
        .O(\rd_data[7]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \rd_data[7]_i_27 
       (.I0(\csr_data_out[11]_i_7_n_0 ),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [7]),
        .O(\rd_data[7]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4545454444444544)) 
    \rd_data[7]_i_28 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\csr_data_out[7]_i_6_n_0 ),
        .I2(\csr_data_out[4]_i_9_n_0 ),
        .I3(\rd_data[7]_i_37_n_0 ),
        .I4(\csr_data_out[30]_i_9_n_0 ),
        .I5(\processor/wb_exception_context[badaddr] [7]),
        .O(\rd_data[7]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[7]_i_29 
       (.I0(\processor/ex_pc [6]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [6]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [6]),
        .O(\rd_data[7]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[7]_i_3 
       (.I0(\rd_data[7]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [7]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[7]_i_8_n_0 ),
        .O(\rd_data[7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \rd_data[7]_i_30 
       (.I0(\processor/mem_exception_context[badaddr] [6]),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .O(\rd_data[7]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000540455555555)) 
    \rd_data[7]_i_31 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\rd_data[7]_i_38_n_0 ),
        .I2(\csr_data_out[30]_i_9_n_0 ),
        .I3(\processor/wb_exception_context[badaddr] [6]),
        .I4(\csr_data_out[4]_i_9_n_0 ),
        .I5(\rd_data[7]_i_39_n_0 ),
        .O(\rd_data[7]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[7]_i_32 
       (.I0(\processor/ex_pc [5]),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/immediate [5]),
        .I3(\processor/execute/alu_x_src [0]),
        .I4(\processor/execute/rs1_forwarded [5]),
        .O(\rd_data[7]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \rd_data[7]_i_33 
       (.I0(\csr_data_out[11]_i_7_n_0 ),
        .I1(\csr_data_out[30]_i_7_n_0 ),
        .I2(\processor/mem_exception_context[badaddr] [5]),
        .O(\rd_data[7]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4545454444444544)) 
    \rd_data[7]_i_34 
       (.I0(\csr_data_out[31]_i_6_n_0 ),
        .I1(\csr_data_out[5]_i_6_n_0 ),
        .I2(\csr_data_out[4]_i_9_n_0 ),
        .I3(\rd_data[7]_i_40_n_0 ),
        .I4(\csr_data_out[30]_i_9_n_0 ),
        .I5(\processor/wb_exception_context[badaddr] [5]),
        .O(\rd_data[7]_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[7]_i_35 
       (.I0(\processor/ex_pc [4]),
        .I1(\processor/execute/shamt [4]),
        .I2(\processor/execute/alu_x_src [1]),
        .I3(\processor/execute/immediate [4]),
        .I4(\processor/execute/alu_x_src [0]),
        .I5(\processor/execute/rs1_forwarded [4]),
        .O(\rd_data[7]_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[7]_i_36 
       (.I0(\processor/ex_pc [7]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [7]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [7]),
        .O(\rd_data[7]_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEAEAEAAA2A2A2AAA)) 
    \rd_data[7]_i_37 
       (.I0(\processor/csr_read_data [7]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded3 ),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/wb_csr_write [0]),
        .I5(\processor/wb_csr_data [7]),
        .O(\rd_data[7]_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEAEAEAAA2A2A2AAA)) 
    \rd_data[7]_i_38 
       (.I0(\processor/csr_read_data [6]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded3 ),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/wb_csr_write [0]),
        .I5(\processor/wb_csr_data [6]),
        .O(\rd_data[7]_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7F7F7FFF)) 
    \rd_data[7]_i_39 
       (.I0(\processor/mem_csr_data [6]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded30_out ),
        .I3(\processor/mem_csr_write [0]),
        .I4(\processor/mem_csr_write [1]),
        .O(\rd_data[7]_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rd_data[7]_i_4 
       (.I0(\rd_data[13]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[9]_i_8_n_0 ),
        .I3(\rd_data[11]_i_9_n_0 ),
        .I4(\rd_data[7]_i_9_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[7]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEAEAEAAA2A2A2AAA)) 
    \rd_data[7]_i_40 
       (.I0(\processor/csr_read_data [5]),
        .I1(\processor/execute/csr_writeable ),
        .I2(\processor/execute/csr_value_forwarded3 ),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/wb_csr_write [0]),
        .I5(\processor/wb_csr_data [5]),
        .O(\rd_data[7]_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rd_data[7]_i_5 
       (.I0(\rd_data[7]_i_10_n_0 ),
        .I1(\processor/execute/alu_y [1]),
        .I2(\rd_data[9]_i_9_n_0 ),
        .O(\rd_data[7]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[7]_i_6 
       (.I0(\rd_data[8]_i_10_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[7]_i_11_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [7]),
        .O(\rd_data[7]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[7]_i_8 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [7]),
        .I3(\processor/execute/alu_y [7]),
        .O(\rd_data[7]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[7]_i_9 
       (.I0(\processor/execute/alu_x [31]),
        .I1(\processor/execute/alu_x [15]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_x [23]),
        .I4(\processor/execute/alu_y [4]),
        .I5(\processor/execute/alu_x [7]),
        .O(\rd_data[7]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[8]_i_1 
       (.I0(\rd_data[8]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[8]_i_3_n_0 ),
        .O(\processor/ex_rd_data [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[8]_i_10 
       (.I0(\rd_data[12]_i_12_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[8]_i_12_n_0 ),
        .I3(\rd_data[14]_i_12_n_0 ),
        .I4(\rd_data[10]_i_13_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[8]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[8]_i_11 
       (.I0(\rd_data[8]_i_13_n_0 ),
        .I1(\csr_data_out[8]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [8]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \rd_data[8]_i_12 
       (.I0(\processor/execute/alu_x [16]),
        .I1(\processor/execute/alu_y [3]),
        .I2(\processor/execute/alu_x [24]),
        .I3(\processor/execute/alu_y [4]),
        .I4(\processor/execute/alu_x [8]),
        .O(\rd_data[8]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[8]_i_13 
       (.I0(\processor/ex_pc [8]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [8]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [8]),
        .O(\rd_data[8]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[8]_i_2 
       (.I0(\rd_data[9]_i_4_n_0 ),
        .I1(\rd_data[8]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[8]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[9]_i_5_n_0 ),
        .O(\rd_data[8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[8]_i_3 
       (.I0(\rd_data[8]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [8]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[8]_i_7_n_0 ),
        .O(\rd_data[8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[8]_i_4 
       (.I0(\rd_data[12]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[8]_i_8_n_0 ),
        .I3(\rd_data[14]_i_8_n_0 ),
        .I4(\rd_data[10]_i_8_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \rd_data[8]_i_5 
       (.I0(\rd_data[10]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[14]_i_9_n_0 ),
        .I3(\rd_data[8]_i_9_n_0 ),
        .I4(\processor/execute/alu_y [1]),
        .O(\rd_data[8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[8]_i_6 
       (.I0(\rd_data[9]_i_10_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[8]_i_10_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [8]),
        .O(\rd_data[8]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[8]_i_7 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [8]),
        .I3(\processor/execute/alu_y [8]),
        .O(\rd_data[8]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[8]_i_8 
       (.I0(\processor/execute/alu_x [31]),
        .I1(\processor/execute/alu_x [16]),
        .I2(\processor/execute/alu_y [3]),
        .I3(\processor/execute/alu_x [24]),
        .I4(\processor/execute/alu_y [4]),
        .I5(\processor/execute/alu_x [8]),
        .O(\rd_data[8]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \rd_data[8]_i_9 
       (.I0(\processor/execute/alu_x [1]),
        .I1(\processor/execute/alu_y [2]),
        .I2(\processor/execute/alu_y [4]),
        .I3(\processor/execute/alu_x [5]),
        .I4(\processor/execute/alu_y [3]),
        .O(\rd_data[8]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \rd_data[9]_i_1 
       (.I0(\rd_data[9]_i_2_n_0 ),
        .I1(\processor/execute/alu_op [2]),
        .I2(\processor/execute/alu_op [1]),
        .I3(\processor/execute/alu_op [3]),
        .I4(\rd_data[9]_i_3_n_0 ),
        .O(\processor/ex_rd_data [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[9]_i_10 
       (.I0(\rd_data[13]_i_12_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[9]_i_12_n_0 ),
        .I3(\rd_data[15]_i_22_n_0 ),
        .I4(\rd_data[11]_i_23_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[9]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30AA30AA3FAA30AA)) 
    \rd_data[9]_i_11 
       (.I0(\rd_data[9]_i_13_n_0 ),
        .I1(\csr_data_out[9]_i_3_n_0 ),
        .I2(\processor/execute/alu_y_src [1]),
        .I3(\processor/execute/alu_y_src [2]),
        .I4(\processor/execute/alu_y_mux/data3 [9]),
        .I5(\processor/execute/alu_y_src [0]),
        .O(\processor/execute/alu_y [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h3300B8B8)) 
    \rd_data[9]_i_12 
       (.I0(\processor/execute/alu_x [25]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [9]),
        .I3(\processor/execute/alu_x [17]),
        .I4(\processor/execute/alu_y [3]),
        .O(\rd_data[9]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \rd_data[9]_i_13 
       (.I0(\processor/ex_pc [9]),
        .I1(\processor/execute/alu_y_src [1]),
        .I2(\processor/execute/immediate [9]),
        .I3(\processor/execute/alu_y_src [0]),
        .I4(\processor/ex_dmem_data_out [9]),
        .O(\rd_data[9]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rd_data[9]_i_2 
       (.I0(\rd_data[10]_i_4_n_0 ),
        .I1(\rd_data[9]_i_4_n_0 ),
        .I2(\rd_data[31]_i_10_n_0 ),
        .I3(\rd_data[9]_i_5_n_0 ),
        .I4(\processor/execute/alu_y [0]),
        .I5(\rd_data[10]_i_5_n_0 ),
        .O(\rd_data[9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888FFFFB8880000)) 
    \rd_data[9]_i_3 
       (.I0(\rd_data[9]_i_6_n_0 ),
        .I1(\processor/execute/alu_op [1]),
        .I2(\processor/execute/alu_op [0]),
        .I3(\processor/execute/alu_instance/data5 [9]),
        .I4(\processor/execute/alu_op [2]),
        .I5(\rd_data[9]_i_7_n_0 ),
        .O(\rd_data[9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[9]_i_4 
       (.I0(\rd_data[13]_i_8_n_0 ),
        .I1(\processor/execute/alu_y [2]),
        .I2(\rd_data[9]_i_8_n_0 ),
        .I3(\rd_data[15]_i_9_n_0 ),
        .I4(\rd_data[11]_i_9_n_0 ),
        .I5(\processor/execute/alu_y [1]),
        .O(\rd_data[9]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rd_data[9]_i_5 
       (.I0(\rd_data[9]_i_9_n_0 ),
        .I1(\processor/execute/alu_y [1]),
        .I2(\rd_data[11]_i_10_n_0 ),
        .O(\rd_data[9]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rd_data[9]_i_6 
       (.I0(\rd_data[10]_i_10_n_0 ),
        .I1(\processor/execute/alu_y [0]),
        .I2(\rd_data[9]_i_10_n_0 ),
        .I3(\processor/execute/alu_op [0]),
        .I4(\processor/execute/alu_instance/data6 [9]),
        .O(\rd_data[9]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5660)) 
    \rd_data[9]_i_7 
       (.I0(\processor/execute/alu_op [1]),
        .I1(\processor/execute/alu_op [0]),
        .I2(\processor/execute/alu_x [9]),
        .I3(\processor/execute/alu_y [9]),
        .O(\rd_data[9]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \rd_data[9]_i_8 
       (.I0(\processor/execute/alu_x [25]),
        .I1(\processor/execute/alu_y [4]),
        .I2(\processor/execute/alu_x [9]),
        .I3(\processor/execute/alu_x [31]),
        .I4(\processor/execute/alu_x [17]),
        .I5(\processor/execute/alu_y [3]),
        .O(\rd_data[9]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \rd_data[9]_i_9 
       (.I0(\processor/execute/alu_x [2]),
        .I1(\processor/execute/alu_y [2]),
        .I2(\processor/execute/alu_y [4]),
        .I3(\processor/execute/alu_x [6]),
        .I4(\processor/execute/alu_y [3]),
        .O(\rd_data[9]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hCCAC)) 
    \rd_data_out[0]_i_1 
       (.I0(\dmem_if/dmem_data_out_reg_n_0_ ),
        .I1(rd_data[0]),
        .I2(\processor/mem_mem_op[1]_repN ),
        .I3(\processor/mem_mem_op [2]),
        .O(\processor/mem_rd_data [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAFCAAAAAA00AAAA)) 
    \rd_data_out[10]_i_1 
       (.I0(rd_data[10]),
        .I1(mem_size[0]),
        .I2(mem_size[1]),
        .I3(\processor/mem_mem_op [2]),
        .I4(\processor/mem_mem_op [1]),
        .I5(\dmem_if/dmem_data_out_reg_n_0_[10] ),
        .O(rd_data_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAFCAAAAAA00AAAA)) 
    \rd_data_out[11]_i_1 
       (.I0(rd_data[11]),
        .I1(mem_size[0]),
        .I2(mem_size[1]),
        .I3(\processor/mem_mem_op [2]),
        .I4(\processor/mem_mem_op [1]),
        .I5(\dmem_if/dmem_data_out_reg_n_0_[11] ),
        .O(\rd_data_out[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAFCAAAAAA00AAAA)) 
    \rd_data_out[12]_i_1 
       (.I0(rd_data[12]),
        .I1(mem_size[0]),
        .I2(mem_size[1]),
        .I3(\processor/mem_mem_op [2]),
        .I4(\processor/mem_mem_op [1]),
        .I5(\dmem_if/dmem_data_out_reg_n_0_[12] ),
        .O(\rd_data_out[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAFCAAAAAA00AAAA)) 
    \rd_data_out[13]_i_1 
       (.I0(rd_data[13]),
        .I1(mem_size[0]),
        .I2(mem_size[1]),
        .I3(\processor/mem_mem_op [2]),
        .I4(\processor/mem_mem_op [1]),
        .I5(\dmem_if/dmem_data_out_reg_n_0_[13] ),
        .O(\rd_data_out[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAFCAAAAAA00AAAA)) 
    \rd_data_out[14]_i_1 
       (.I0(rd_data[14]),
        .I1(mem_size[0]),
        .I2(mem_size[1]),
        .I3(\processor/mem_mem_op [2]),
        .I4(\processor/mem_mem_op [1]),
        .I5(\dmem_if/dmem_data_out_reg_n_0_[14] ),
        .O(\rd_data_out[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \rd_data_out[15]_i_1 
       (.I0(\rd_data_out[15]_i_3_n_0 ),
        .I1(reset),
        .O(\rd_data_out[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAFCAAAAAA00AAAA)) 
    \rd_data_out[15]_i_2 
       (.I0(rd_data[15]),
        .I1(mem_size[0]),
        .I2(mem_size[1]),
        .I3(\processor/mem_mem_op [2]),
        .I4(\processor/mem_mem_op [1]),
        .I5(p_1_in0),
        .O(\rd_data_out[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFEFFFFFFFFF)) 
    \rd_data_out[15]_i_3 
       (.I0(\mem_size[0]_repN ),
        .I1(\mem_size[1]_repN ),
        .I2(\processor/mem_mem_op[1]_repN ),
        .I3(\processor/mem_mem_op [0]),
        .I4(\processor/mem_mem_op [2]),
        .I5(p_0_in0_repN),
        .O(\rd_data_out[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000F333AAAAAAAA)) 
    \rd_data_out[16]_i_1 
       (.I0(rd_data[16]),
        .I1(\rd_data_out[31]_i_2_n_0 ),
        .I2(\dmem_if/dmem_data_out_reg_n_0_[16] ),
        .I3(mem_size[1]),
        .I4(\rd_data_out[31]_i_3_n_0 ),
        .I5(\rd_data_out[31]_i_4_n_0 ),
        .O(\processor/mem_rd_data [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000F333AAAAAAAA)) 
    \rd_data_out[17]_i_1 
       (.I0(rd_data[17]),
        .I1(\rd_data_out[31]_i_2_n_0_repN ),
        .I2(\dmem_if/dmem_data_out_reg_n_0_[17] ),
        .I3(\mem_size[1]_repN ),
        .I4(\rd_data_out[31]_i_3_n_0 ),
        .I5(\rd_data_out[31]_i_4_n_0 ),
        .O(\processor/mem_rd_data [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000F333AAAAAAAA)) 
    \rd_data_out[18]_i_1 
       (.I0(rd_data[18]),
        .I1(\rd_data_out[31]_i_2_n_0_repN ),
        .I2(\dmem_if/dmem_data_out_reg_n_0_[18] ),
        .I3(\mem_size[1]_repN ),
        .I4(\rd_data_out[31]_i_3_n_0 ),
        .I5(\rd_data_out[31]_i_4_n_0 ),
        .O(\processor/mem_rd_data [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000F333AAAAAAAA)) 
    \rd_data_out[19]_i_1 
       (.I0(rd_data[19]),
        .I1(\rd_data_out[31]_i_2_n_0_repN ),
        .I2(\dmem_if/dmem_data_out_reg_n_0_[19] ),
        .I3(\mem_size[1]_repN ),
        .I4(\rd_data_out[31]_i_3_n_0 ),
        .I5(\rd_data_out[31]_i_4_n_0 ),
        .O(\processor/mem_rd_data [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hCCAC)) 
    \rd_data_out[1]_i_1 
       (.I0(\dmem_if/dmem_data_out_reg_n_0_[1] ),
        .I1(rd_data[1]),
        .I2(\processor/mem_mem_op[1]_repN ),
        .I3(\processor/mem_mem_op [2]),
        .O(\processor/mem_rd_data [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000F333AAAAAAAA)) 
    \rd_data_out[20]_i_1 
       (.I0(rd_data[20]),
        .I1(\rd_data_out[31]_i_2_n_0 ),
        .I2(\dmem_if/dmem_data_out_reg_n_0_[20] ),
        .I3(\mem_size[1]_repN_1 ),
        .I4(\rd_data_out[31]_i_3_n_0 ),
        .I5(\rd_data_out[31]_i_4_n_0 ),
        .O(\processor/mem_rd_data [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000F333AAAAAAAA)) 
    \rd_data_out[21]_i_1 
       (.I0(rd_data[21]),
        .I1(\rd_data_out[31]_i_2_n_0_repN ),
        .I2(\dmem_if/dmem_data_out_reg_n_0_[21] ),
        .I3(\mem_size[1]_repN ),
        .I4(\rd_data_out[31]_i_3_n_0 ),
        .I5(\rd_data_out[31]_i_4_n_0 ),
        .O(\processor/mem_rd_data [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000F333AAAAAAAA)) 
    \rd_data_out[22]_i_1 
       (.I0(rd_data[22]),
        .I1(\rd_data_out[31]_i_2_n_0 ),
        .I2(\dmem_if/dmem_data_out_reg_n_0_[22] ),
        .I3(\mem_size[1]_repN ),
        .I4(\rd_data_out[31]_i_3_n_0 ),
        .I5(\rd_data_out[31]_i_4_n_0 ),
        .O(\processor/mem_rd_data [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000F333AAAAAAAA)) 
    \rd_data_out[23]_i_1 
       (.I0(rd_data[23]),
        .I1(\rd_data_out[31]_i_2_n_0_repN ),
        .I2(\dmem_if/dmem_data_out_reg_n_0_[23] ),
        .I3(\mem_size[1]_repN ),
        .I4(\rd_data_out[31]_i_3_n_0 ),
        .I5(\rd_data_out[31]_i_4_n_0 ),
        .O(\processor/mem_rd_data [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000F333AAAAAAAA)) 
    \rd_data_out[24]_i_1 
       (.I0(rd_data[24]),
        .I1(\rd_data_out[31]_i_2_n_0_repN ),
        .I2(\dmem_if/dmem_data_out_reg_n_0_[24] ),
        .I3(\mem_size[1]_repN ),
        .I4(\rd_data_out[31]_i_3_n_0 ),
        .I5(\rd_data_out[31]_i_4_n_0 ),
        .O(\processor/mem_rd_data [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000F333AAAAAAAA)) 
    \rd_data_out[25]_i_1 
       (.I0(rd_data[25]),
        .I1(\rd_data_out[31]_i_2_n_0 ),
        .I2(\dmem_if/dmem_data_out_reg_n_0_[25] ),
        .I3(\mem_size[1]_repN ),
        .I4(\rd_data_out[31]_i_3_n_0 ),
        .I5(\rd_data_out[31]_i_4_n_0 ),
        .O(\processor/mem_rd_data [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000F333AAAAAAAA)) 
    \rd_data_out[26]_i_1 
       (.I0(rd_data[26]),
        .I1(\rd_data_out[31]_i_2_n_0 ),
        .I2(\dmem_if/dmem_data_out_reg_n_0_[26] ),
        .I3(\mem_size[1]_repN_1 ),
        .I4(\rd_data_out[31]_i_3_n_0 ),
        .I5(\rd_data_out[31]_i_4_n_0 ),
        .O(\processor/mem_rd_data [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000F333AAAAAAAA)) 
    \rd_data_out[27]_i_1 
       (.I0(rd_data[27]),
        .I1(\rd_data_out[31]_i_2_n_0 ),
        .I2(\dmem_if/dmem_data_out_reg_n_0_[27] ),
        .I3(\mem_size[1]_repN_1 ),
        .I4(\rd_data_out[31]_i_3_n_0 ),
        .I5(\rd_data_out[31]_i_4_n_0 ),
        .O(\processor/mem_rd_data [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000F333AAAAAAAA)) 
    \rd_data_out[28]_i_1 
       (.I0(rd_data[28]),
        .I1(\rd_data_out[31]_i_2_n_0 ),
        .I2(\dmem_if/dmem_data_out_reg_n_0_[28] ),
        .I3(\mem_size[1]_repN_1 ),
        .I4(\rd_data_out[31]_i_3_n_0 ),
        .I5(\rd_data_out[31]_i_4_n_0 ),
        .O(\processor/mem_rd_data [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000F333AAAAAAAA)) 
    \rd_data_out[29]_i_1 
       (.I0(rd_data[29]),
        .I1(\rd_data_out[31]_i_2_n_0 ),
        .I2(\dmem_if/dmem_data_out_reg_n_0_[29] ),
        .I3(\mem_size[1]_repN ),
        .I4(\rd_data_out[31]_i_3_n_0 ),
        .I5(\rd_data_out[31]_i_4_n_0 ),
        .O(\processor/mem_rd_data [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hCCAC)) 
    \rd_data_out[2]_i_1 
       (.I0(\dmem_if/dmem_data_out_reg_n_0_[2] ),
        .I1(rd_data[2]),
        .I2(\processor/mem_mem_op[1]_repN ),
        .I3(\processor/mem_mem_op [2]),
        .O(\processor/mem_rd_data [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000F333AAAAAAAA)) 
    \rd_data_out[30]_i_1 
       (.I0(rd_data[30]),
        .I1(\rd_data_out[31]_i_2_n_0 ),
        .I2(\dmem_if/dmem_data_out_reg_n_0_[30] ),
        .I3(\mem_size[1]_repN ),
        .I4(\rd_data_out[31]_i_3_n_0 ),
        .I5(\rd_data_out[31]_i_4_n_0 ),
        .O(\processor/mem_rd_data [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000F333AAAAAAAA)) 
    \rd_data_out[31]_i_1 
       (.I0(rd_data[31]),
        .I1(\rd_data_out[31]_i_2_n_0 ),
        .I2(\dmem_if/dmem_data_out_reg_n_0_[31] ),
        .I3(\mem_size[1]_repN ),
        .I4(\rd_data_out[31]_i_3_n_0 ),
        .I5(\rd_data_out[31]_i_4_n_0 ),
        .O(\processor/mem_rd_data [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    \rd_data_out[31]_i_2 
       (.I0(mem_size[1]),
        .I1(\processor/mem_mem_op [2]),
        .I2(\processor/mem_mem_op [0]),
        .I3(\processor/mem_mem_op[1]_repN ),
        .O(\rd_data_out[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "rd_data_out[31]_i_2" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    \rd_data_out[31]_i_2_replica 
       (.I0(\mem_size[1]_repN_2 ),
        .I1(\processor/mem_mem_op [2]),
        .I2(\processor/mem_mem_op [0]),
        .I3(\processor/mem_mem_op[1]_repN ),
        .O(\rd_data_out[31]_i_2_n_0_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h001D)) 
    \rd_data_out[31]_i_3 
       (.I0(p_0_in0_repN),
        .I1(mem_size[0]),
        .I2(p_1_in0),
        .I3(mem_size[1]),
        .O(\rd_data_out[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \rd_data_out[31]_i_4 
       (.I0(\processor/mem_mem_op[1]_repN ),
        .I1(\processor/mem_mem_op [2]),
        .O(\rd_data_out[31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hCCAC)) 
    \rd_data_out[3]_i_1 
       (.I0(\dmem_if/dmem_data_out_reg_n_0_[3] ),
        .I1(rd_data[3]),
        .I2(\processor/mem_mem_op[1]_repN_1 ),
        .I3(\processor/mem_mem_op [2]),
        .O(\processor/mem_rd_data [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hCCAC)) 
    \rd_data_out[4]_i_1 
       (.I0(\dmem_if/dmem_data_out_reg_n_0_[4] ),
        .I1(rd_data[4]),
        .I2(\processor/mem_mem_op[1]_repN_1 ),
        .I3(\processor/mem_mem_op [2]),
        .O(\processor/mem_rd_data [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hCCAC)) 
    \rd_data_out[5]_i_1 
       (.I0(\dmem_if/dmem_data_out_reg_n_0_[5] ),
        .I1(rd_data[5]),
        .I2(\processor/mem_mem_op[1]_repN_2 ),
        .I3(\processor/mem_mem_op [2]),
        .O(\processor/mem_rd_data [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hCCAC)) 
    \rd_data_out[6]_i_1 
       (.I0(\dmem_if/dmem_data_out_reg_n_0_[6] ),
        .I1(rd_data[6]),
        .I2(\processor/mem_mem_op[1]_repN_1 ),
        .I3(\processor/mem_mem_op [2]),
        .O(\processor/mem_rd_data [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hCCAC)) 
    \rd_data_out[7]_i_1 
       (.I0(p_0_in0),
        .I1(rd_data[7]),
        .I2(\processor/mem_mem_op[1]_repN ),
        .I3(\processor/mem_mem_op [2]),
        .O(\processor/mem_rd_data [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "rd_data_out[7]_i_1" *) 
  LUT4 #(
    .INIT(16'hCCAC)) 
    \rd_data_out[7]_i_1_replica 
       (.I0(p_0_in0),
        .I1(rd_data[7]),
        .I2(\processor/mem_mem_op[1]_repN ),
        .I3(\processor/mem_mem_op [2]),
        .O(\processor/mem_rd_data[7]_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "rd_data_out[7]_i_1" *) 
  LUT4 #(
    .INIT(16'hCCAC)) 
    \rd_data_out[7]_i_1_replica_1 
       (.I0(p_0_in0),
        .I1(rd_data[7]),
        .I2(\processor/mem_mem_op[1]_repN ),
        .I3(\processor/mem_mem_op [2]),
        .O(\processor/mem_rd_data[7]_repN_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAFCAAAAAA00AAAA)) 
    \rd_data_out[8]_i_1 
       (.I0(rd_data[8]),
        .I1(mem_size[0]),
        .I2(mem_size[1]),
        .I3(\processor/mem_mem_op [2]),
        .I4(\processor/mem_mem_op [1]),
        .I5(\dmem_if/dmem_data_out_reg_n_0_[8] ),
        .O(\rd_data_out[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAFCAAAAAA00AAAA)) 
    \rd_data_out[9]_i_1 
       (.I0(rd_data[9]),
        .I1(mem_size[0]),
        .I2(mem_size[1]),
        .I3(\processor/mem_mem_op [2]),
        .I4(\processor/mem_mem_op [1]),
        .I5(\dmem_if/dmem_data_out_reg_n_0_[9] ),
        .O(\rd_data_out[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \rd_data_reg[0]_i_1 
       (.I0(\rd_data[0]_i_2_n_0 ),
        .I1(\rd_data[0]_i_3_n_0 ),
        .O(\processor/ex_rd_data [0]),
        .S(\processor/execute/alu_op [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[0]_i_10 
       (.CI(\rd_data_reg[0]_i_22_n_0 ),
        .CO({\processor/execute/alu_instance/data3 ,\rd_data_reg[0]_i_10_n_1 ,\rd_data_reg[0]_i_10_n_2 ,\rd_data_reg[0]_i_10_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\rd_data[0]_i_23_n_0 ,\rd_data[0]_i_15_n_0 ,\rd_data[0]_i_16_n_0 ,\rd_data[0]_i_17_n_0 }),
        .S({\rd_data[0]_i_24_n_0 ,\rd_data[0]_i_25_n_0 ,\rd_data[0]_i_26_n_0 ,\rd_data[0]_i_27_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[0]_i_13 
       (.CI(\rd_data_reg[0]_i_30_n_0 ),
        .CO(rd_data_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\rd_data[0]_i_31_n_0 ,\rd_data[0]_i_32_n_0 ,\rd_data[0]_i_33_n_0 ,\rd_data[0]_i_34_n_0 }),
        .S({\rd_data[0]_i_35_n_0 ,\rd_data[0]_i_36_n_0 ,\rd_data[0]_i_37_n_0 ,\rd_data[0]_i_38_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[0]_i_22 
       (.CI(\rd_data_reg[0]_i_39_n_0 ),
        .CO({\rd_data_reg[0]_i_22_n_0 ,\rd_data_reg[0]_i_22_n_1 ,\rd_data_reg[0]_i_22_n_2 ,\rd_data_reg[0]_i_22_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\rd_data[0]_i_31_n_0 ,\rd_data[0]_i_32_n_0 ,\rd_data[0]_i_33_n_0 ,\rd_data[0]_i_34_n_0 }),
        .S({\rd_data[0]_i_40_n_0 ,\rd_data[0]_i_41_n_0 ,\rd_data[0]_i_42_n_0 ,\rd_data[0]_i_43_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[0]_i_30 
       (.CI(\rd_data_reg[0]_i_44_n_0 ),
        .CO({\rd_data_reg[0]_i_30_n_0 ,\rd_data_reg[0]_i_30_n_1 ,\rd_data_reg[0]_i_30_n_2 ,\rd_data_reg[0]_i_30_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\rd_data[0]_i_45_n_0 ,\rd_data[0]_i_46_n_0 ,\rd_data[0]_i_47_n_0 ,\rd_data[0]_i_48_n_0 }),
        .S({\rd_data[0]_i_49_n_0 ,\rd_data[0]_i_50_n_0 ,\rd_data[0]_i_51_n_0 ,\rd_data[0]_i_52_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[0]_i_39 
       (.CI(\rd_data_reg[0]_i_53_n_0 ),
        .CO({\rd_data_reg[0]_i_39_n_0 ,\rd_data_reg[0]_i_39_n_1 ,\rd_data_reg[0]_i_39_n_2 ,\rd_data_reg[0]_i_39_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\rd_data[0]_i_45_n_0 ,\rd_data[0]_i_46_n_0 ,\rd_data[0]_i_47_n_0 ,\rd_data[0]_i_48_n_0 }),
        .S({\rd_data[0]_i_54_n_0 ,\rd_data[0]_i_55_n_0 ,\rd_data[0]_i_56_n_0 ,\rd_data[0]_i_57_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[0]_i_44 
       (.CI(\<const0>__0__0 ),
        .CO({\rd_data_reg[0]_i_44_n_0 ,\rd_data_reg[0]_i_44_n_1 ,\rd_data_reg[0]_i_44_n_2 ,\rd_data_reg[0]_i_44_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\rd_data[0]_i_58_n_0 ,\rd_data[0]_i_59_n_0 ,\rd_data[0]_i_60_n_0 ,\rd_data[0]_i_61_n_0 }),
        .S({\rd_data[0]_i_62_n_0 ,\rd_data[0]_i_63_n_0 ,\rd_data[0]_i_64_n_0 ,\rd_data[0]_i_65_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[0]_i_53 
       (.CI(\<const0>__0__0 ),
        .CO({\rd_data_reg[0]_i_53_n_0 ,\rd_data_reg[0]_i_53_n_1 ,\rd_data_reg[0]_i_53_n_2 ,\rd_data_reg[0]_i_53_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\rd_data[0]_i_58_n_0 ,\rd_data[0]_i_59_n_0 ,\rd_data[0]_i_60_n_0 ,\rd_data[0]_i_61_n_0 }),
        .S({\rd_data[0]_i_66_n_0 ,\rd_data[0]_i_67_n_0 ,\rd_data[0]_i_68_n_0 ,\rd_data[0]_i_69_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[0]_i_9 
       (.CI(rd_data_reg[3]),
        .CO({\processor/execute/alu_instance/data4 ,\rd_data_reg[0]_i_9_n_1 ,\rd_data_reg[0]_i_9_n_2 ,\rd_data_reg[0]_i_9_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\rd_data[0]_i_14_n_0 ,\rd_data[0]_i_15_n_0 ,\rd_data[0]_i_16_n_0 ,\rd_data[0]_i_17_n_0 }),
        .S({\rd_data[0]_i_18_n_0 ,\rd_data[0]_i_19_n_0 ,\rd_data[0]_i_20_n_0 ,\rd_data[0]_i_21_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[11]_i_12 
       (.CI(\rd_data_reg[7]_i_12_n_0 ),
        .CO({\rd_data_reg[11]_i_12_n_0 ,\rd_data_reg[11]_i_12_n_1 ,\rd_data_reg[11]_i_12_n_2 ,\rd_data_reg[11]_i_12_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\processor/execute/alu_x [11:8]),
        .O(\processor/execute/alu_instance/data6 [11:8]),
        .S({\rd_data[11]_i_24_n_0 ,\rd_data[11]_i_25_n_0 ,\rd_data[11]_i_26_n_0 ,\rd_data[11]_i_27_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[11]_i_40 
       (.CI(\rd_data_reg[2]_i_11_n_0 ),
        .CO({\rd_data_reg[11]_i_40_n_0 ,\rd_data_reg[11]_i_40_n_1 ,\rd_data_reg[11]_i_40_n_2 ,\rd_data_reg[11]_i_40_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\processor/execute/alu_x_mux/data3 [8:5]),
        .S(\processor/ex_pc [8:5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[11]_i_7 
       (.CI(\rd_data_reg[7]_i_7_n_0 ),
        .CO({\rd_data_reg[11]_i_7_n_0 ,\rd_data_reg[11]_i_7_n_1 ,\rd_data_reg[11]_i_7_n_2 ,\rd_data_reg[11]_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\processor/execute/alu_x [11:8]),
        .O(\processor/execute/alu_instance/data5 [11:8]),
        .S({\rd_data[11]_i_17_n_0 ,\rd_data[11]_i_18_n_0 ,\rd_data[11]_i_19_n_0 ,\rd_data[11]_i_20_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[12]_i_14 
       (.CI(\rd_data_reg[8]_i_14_n_0 ),
        .CO({\rd_data_reg[12]_i_14_n_0 ,\rd_data_reg[12]_i_14_n_1 ,\rd_data_reg[12]_i_14_n_2 ,\rd_data_reg[12]_i_14_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\processor/execute/alu_y_mux/data3 [12:9]),
        .S(\processor/ex_pc [12:9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[15]_i_12 
       (.CI(\rd_data_reg[11]_i_12_n_0 ),
        .CO({\rd_data_reg[15]_i_12_n_0 ,\rd_data_reg[15]_i_12_n_1 ,\rd_data_reg[15]_i_12_n_2 ,\rd_data_reg[15]_i_12_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\processor/execute/alu_x [15:12]),
        .O(\processor/execute/alu_instance/data6 [15:12]),
        .S({\rd_data[15]_i_23_n_0 ,\rd_data[15]_i_24_n_0 ,\rd_data[15]_i_25_n_0 ,\rd_data[15]_i_26_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[15]_i_39 
       (.CI(\rd_data_reg[11]_i_40_n_0 ),
        .CO({\rd_data_reg[15]_i_39_n_0 ,\rd_data_reg[15]_i_39_n_1 ,\rd_data_reg[15]_i_39_n_2 ,\rd_data_reg[15]_i_39_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\processor/execute/alu_x_mux/data3 [12:9]),
        .S(\processor/ex_pc [12:9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[15]_i_7 
       (.CI(\rd_data_reg[11]_i_7_n_0 ),
        .CO({\rd_data_reg[15]_i_7_n_0 ,\rd_data_reg[15]_i_7_n_1 ,\rd_data_reg[15]_i_7_n_2 ,\rd_data_reg[15]_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\processor/execute/alu_x [15:12]),
        .O(\processor/execute/alu_instance/data5 [15:12]),
        .S({\rd_data[15]_i_17_n_0 ,\rd_data[15]_i_18_n_0 ,\rd_data[15]_i_19_n_0 ,\rd_data[15]_i_20_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[16]_i_15 
       (.CI(\rd_data_reg[12]_i_14_n_0 ),
        .CO({\rd_data_reg[16]_i_15_n_0 ,\rd_data_reg[16]_i_15_n_1 ,\rd_data_reg[16]_i_15_n_2 ,\rd_data_reg[16]_i_15_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\processor/execute/alu_y_mux/data3 [16:13]),
        .S(\processor/ex_pc [16:13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[19]_i_13 
       (.CI(\rd_data_reg[15]_i_12_n_0 ),
        .CO({\rd_data_reg[19]_i_13_n_0 ,\rd_data_reg[19]_i_13_n_1 ,\rd_data_reg[19]_i_13_n_2 ,\rd_data_reg[19]_i_13_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\processor/execute/alu_x [19:16]),
        .O(\processor/execute/alu_instance/data6 [19:16]),
        .S({\rd_data[19]_i_25_n_0 ,\rd_data[19]_i_26_n_0 ,\rd_data[19]_i_27_n_0 ,\rd_data[19]_i_28_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[19]_i_41 
       (.CI(\rd_data_reg[15]_i_39_n_0 ),
        .CO({\rd_data_reg[19]_i_41_n_0 ,\rd_data_reg[19]_i_41_n_1 ,\rd_data_reg[19]_i_41_n_2 ,\rd_data_reg[19]_i_41_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\processor/execute/alu_x_mux/data3 [16:13]),
        .S(\processor/ex_pc [16:13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[19]_i_7 
       (.CI(\rd_data_reg[15]_i_7_n_0 ),
        .CO({\rd_data_reg[19]_i_7_n_0 ,\rd_data_reg[19]_i_7_n_1 ,\rd_data_reg[19]_i_7_n_2 ,\rd_data_reg[19]_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\processor/execute/alu_x [19:16]),
        .O(\processor/execute/alu_instance/data5 [19:16]),
        .S({\rd_data[19]_i_18_n_0 ,\rd_data[19]_i_19_n_0 ,\rd_data[19]_i_20_n_0 ,\rd_data[19]_i_21_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \rd_data_reg[1]_i_1 
       (.I0(\rd_data[1]_i_2_n_0 ),
        .I1(\rd_data[1]_i_3_n_0 ),
        .O(\processor/ex_rd_data [1]),
        .S(\processor/execute/alu_op [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[20]_i_15 
       (.CI(\rd_data_reg[16]_i_15_n_0 ),
        .CO({\rd_data_reg[20]_i_15_n_0 ,\rd_data_reg[20]_i_15_n_1 ,\rd_data_reg[20]_i_15_n_2 ,\rd_data_reg[20]_i_15_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\processor/execute/alu_y_mux/data3 [20:17]),
        .S(\processor/ex_pc [20:17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[23]_i_12 
       (.CI(\rd_data_reg[19]_i_13_n_0 ),
        .CO({\rd_data_reg[23]_i_12_n_0 ,\rd_data_reg[23]_i_12_n_1 ,\rd_data_reg[23]_i_12_n_2 ,\rd_data_reg[23]_i_12_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\processor/execute/alu_x [23:20]),
        .O(\processor/execute/alu_instance/data6 [23:20]),
        .S({\rd_data[23]_i_23_n_0 ,\rd_data[23]_i_24_n_0 ,\rd_data[23]_i_25_n_0 ,\rd_data[23]_i_26_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[23]_i_39 
       (.CI(\rd_data_reg[19]_i_41_n_0 ),
        .CO({\rd_data_reg[23]_i_39_n_0 ,\rd_data_reg[23]_i_39_n_1 ,\rd_data_reg[23]_i_39_n_2 ,\rd_data_reg[23]_i_39_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\processor/execute/alu_x_mux/data3 [20:17]),
        .S(\processor/ex_pc [20:17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[23]_i_7 
       (.CI(\rd_data_reg[19]_i_7_n_0 ),
        .CO({\rd_data_reg[23]_i_7_n_0 ,\rd_data_reg[23]_i_7_n_1 ,\rd_data_reg[23]_i_7_n_2 ,\rd_data_reg[23]_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\processor/execute/alu_x [23:20]),
        .O(\processor/execute/alu_instance/data5 [23:20]),
        .S({\rd_data[23]_i_17_n_0 ,\rd_data[23]_i_18_n_0 ,\rd_data[23]_i_19_n_0 ,\rd_data[23]_i_20_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[24]_i_14 
       (.CI(\rd_data_reg[20]_i_15_n_0 ),
        .CO({\rd_data_reg[24]_i_14_n_0 ,\rd_data_reg[24]_i_14_n_1 ,\rd_data_reg[24]_i_14_n_2 ,\rd_data_reg[24]_i_14_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\processor/execute/alu_y_mux/data3 [24:21]),
        .S(\processor/ex_pc [24:21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[27]_i_13 
       (.CI(\rd_data_reg[23]_i_12_n_0 ),
        .CO({\rd_data_reg[27]_i_13_n_0 ,\rd_data_reg[27]_i_13_n_1 ,\rd_data_reg[27]_i_13_n_2 ,\rd_data_reg[27]_i_13_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\processor/execute/alu_x [27:24]),
        .O(\processor/execute/alu_instance/data6 [27:24]),
        .S({\rd_data[27]_i_24_n_0 ,\rd_data[27]_i_25_n_0 ,\rd_data[27]_i_26_n_0 ,\rd_data[27]_i_27_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[27]_i_40 
       (.CI(\rd_data_reg[23]_i_39_n_0 ),
        .CO({\rd_data_reg[27]_i_40_n_0 ,\rd_data_reg[27]_i_40_n_1 ,\rd_data_reg[27]_i_40_n_2 ,\rd_data_reg[27]_i_40_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\processor/execute/alu_x_mux/data3 [24:21]),
        .S(\processor/ex_pc [24:21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[27]_i_7 
       (.CI(\rd_data_reg[23]_i_7_n_0 ),
        .CO({\rd_data_reg[27]_i_7_n_0 ,\rd_data_reg[27]_i_7_n_1 ,\rd_data_reg[27]_i_7_n_2 ,\rd_data_reg[27]_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\processor/execute/alu_x [27:24]),
        .O(\processor/execute/alu_instance/data5 [27:24]),
        .S({\rd_data[27]_i_18_n_0 ,\rd_data[27]_i_19_n_0 ,\rd_data[27]_i_20_n_0 ,\rd_data[27]_i_21_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \rd_data_reg[2]_i_1 
       (.I0(\rd_data[2]_i_2_n_0 ),
        .I1(\rd_data[2]_i_3_n_0 ),
        .O(\processor/ex_rd_data [2]),
        .S(\processor/execute/alu_op [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[2]_i_11 
       (.CI(\<const0>__0__0 ),
        .CO({\rd_data_reg[2]_i_11_n_0 ,\rd_data_reg[2]_i_11_n_1 ,\rd_data_reg[2]_i_11_n_2 ,\rd_data_reg[2]_i_11_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\processor/ex_pc [2],\<const0>__0__0 }),
        .O(\processor/execute/alu_x_mux/data3 [4:1]),
        .S({\processor/ex_pc [4:3],\rd_data[2]_i_17_n_0 ,\processor/ex_pc [1]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[2]_i_13 
       (.CI(\<const0>__0__0 ),
        .CO({\rd_data_reg[2]_i_13_n_0 ,\rd_data_reg[2]_i_13_n_1 ,\rd_data_reg[2]_i_13_n_2 ,\rd_data_reg[2]_i_13_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\processor/ex_pc [2],\<const0>__0__0 }),
        .O(\processor/execute/alu_y_mux/data3 [4:1]),
        .S({\processor/ex_pc [4:3],\rd_data[2]_i_21_n_0 ,\processor/ex_pc [1]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[30]_i_7 
       (.CI(\rd_data_reg[27]_i_7_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\processor/execute/alu_x [30:28]}),
        .O(\processor/execute/alu_instance/data5 [31:28]),
        .S({\rd_data[30]_i_16_n_0 ,\rd_data[30]_i_17_n_0 ,\rd_data[30]_i_18_n_0 ,\rd_data[30]_i_19_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \rd_data_reg[31]_i_1 
       (.I0(\rd_data[31]_i_2_n_0 ),
        .I1(\rd_data[31]_i_3_n_0 ),
        .O(\processor/ex_rd_data [31]),
        .S(\processor/execute/alu_op [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[31]_i_13 
       (.CI(\rd_data_reg[27]_i_13_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\processor/execute/alu_x [30:28]}),
        .O(\processor/execute/alu_instance/data6 [31:28]),
        .S({\rd_data[31]_i_28_n_0 ,\rd_data[31]_i_29_n_0 ,\rd_data[31]_i_30_n_0 ,\rd_data[31]_i_31_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[31]_i_15 
       (.CI(\rd_data_reg[31]_i_32_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\rd_data_reg[31]_i_15_n_4 ,\processor/execute/alu_x_mux/data3 [31:29]}),
        .S({\<const0>__0__0 ,\processor/ex_pc [31:29]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[31]_i_17 
       (.CI(\rd_data_reg[31]_i_36_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\rd_data_reg[31]_i_17_n_4 ,\processor/execute/alu_y_mux/data3 [31:29]}),
        .S({\<const0>__0__0 ,\processor/ex_pc [31:29]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[31]_i_32 
       (.CI(\rd_data_reg[27]_i_40_n_0 ),
        .CO({\rd_data_reg[31]_i_32_n_0 ,\rd_data_reg[31]_i_32_n_1 ,\rd_data_reg[31]_i_32_n_2 ,\rd_data_reg[31]_i_32_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\processor/execute/alu_x_mux/data3 [28:25]),
        .S(\processor/ex_pc [28:25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[31]_i_36 
       (.CI(\rd_data_reg[24]_i_14_n_0 ),
        .CO({\rd_data_reg[31]_i_36_n_0 ,\rd_data_reg[31]_i_36_n_1 ,\rd_data_reg[31]_i_36_n_2 ,\rd_data_reg[31]_i_36_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\processor/execute/alu_y_mux/data3 [28:25]),
        .S(\processor/ex_pc [28:25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[3]_i_12 
       (.CI(\<const0>__0__0 ),
        .CO({\rd_data_reg[3]_i_12_n_0 ,\rd_data_reg[3]_i_12_n_1 ,\rd_data_reg[3]_i_12_n_2 ,\rd_data_reg[3]_i_12_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI(\processor/execute/alu_x [3:0]),
        .O(\processor/execute/alu_instance/data6 [3:0]),
        .S({\rd_data[3]_i_21_n_0 ,\rd_data[3]_i_22_n_0 ,\rd_data[3]_i_23_n_0 ,\rd_data[3]_i_24_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[3]_i_7 
       (.CI(\<const0>__0__0 ),
        .CO({\rd_data_reg[3]_i_7_n_0 ,\rd_data_reg[3]_i_7_n_1 ,\rd_data_reg[3]_i_7_n_2 ,\rd_data_reg[3]_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\processor/execute/alu_x [3:0]),
        .O(\processor/execute/alu_instance/data5 [3:0]),
        .S({\rd_data[3]_i_14_n_0 ,\rd_data[3]_i_15_n_0 ,\rd_data[3]_i_16_n_0 ,\rd_data[3]_i_17_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[7]_i_12 
       (.CI(\rd_data_reg[3]_i_12_n_0 ),
        .CO({\rd_data_reg[7]_i_12_n_0 ,\rd_data_reg[7]_i_12_n_1 ,\rd_data_reg[7]_i_12_n_2 ,\rd_data_reg[7]_i_12_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\processor/execute/alu_x [7:4]),
        .O(\processor/execute/alu_instance/data6 [7:4]),
        .S({\rd_data[7]_i_22_n_0 ,\rd_data[7]_i_23_n_0 ,\rd_data[7]_i_24_n_0 ,\rd_data[7]_i_25_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[7]_i_7 
       (.CI(\rd_data_reg[3]_i_7_n_0 ),
        .CO({\rd_data_reg[7]_i_7_n_0 ,\rd_data_reg[7]_i_7_n_1 ,\rd_data_reg[7]_i_7_n_2 ,\rd_data_reg[7]_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\processor/execute/alu_x [7:4]),
        .O(\processor/execute/alu_instance/data5 [7:4]),
        .S({\rd_data[7]_i_17_n_0 ,\rd_data[7]_i_18_n_0 ,\rd_data[7]_i_19_n_0 ,\rd_data[7]_i_20_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rd_data_reg[8]_i_14 
       (.CI(\rd_data_reg[2]_i_13_n_0 ),
        .CO({\rd_data_reg[8]_i_14_n_0 ,\rd_data_reg[8]_i_14_n_1 ,\rd_data_reg[8]_i_14_n_2 ,\rd_data_reg[8]_i_14_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\processor/execute/alu_y_mux/data3 [8:5]),
        .S(\processor/ex_pc [8:5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00CC0F0008000F03)) 
    rd_write_out_i_1
       (.I0(rd_write_out_i_2_n_0),
        .I1(\processor/decode/instruction_reg_n_0_[5] ),
        .I2(\processor/decode/instruction_reg_n_0_[3] ),
        .I3(\processor/decode/instruction_reg_n_0_[4] ),
        .I4(\processor/decode/instruction_reg_n_0_[6] ),
        .I5(\processor/decode/instruction_reg_n_0_ ),
        .O(\processor/id_rd_write ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    rd_write_out_i_2
       (.I0(\processor/id_csr_use_immediate ),
        .I1(\processor/decode/instruction_reg_n_0_ ),
        .I2(\processor/id_funct3 [0]),
        .I3(\processor/id_funct3 [1]),
        .O(rd_write_out_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFA0008)) 
    read_ack_i_1
       (.I0(\icache/state_reg_n_0_[1] ),
        .I1(icache_inputs),
        .I2(\icache/state_reg_n_0_ ),
        .I3(\icache/state_reg_n_0_[2] ),
        .I4(\icache/read_ack ),
        .O(read_ack_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    read_data_out2_carry_i_1
       (.I0(\processor/wb_csr_address [9]),
        .I1(\csr_addr[9]_i_1_n_0 ),
        .I2(\csr_addr[11]_i_1_n_0 ),
        .I3(\processor/wb_csr_address [11]),
        .I4(\csr_addr[10]_i_1_n_0 ),
        .I5(\processor/wb_csr_address [10]),
        .O(read_data_out2_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    read_data_out2_carry_i_2
       (.I0(\processor/wb_csr_address [6]),
        .I1(\csr_addr[6]_i_1_n_0 ),
        .I2(\csr_addr[8]_i_1_n_0 ),
        .I3(\processor/wb_csr_address [8]),
        .I4(\csr_addr[7]_i_1_n_0 ),
        .I5(\processor/wb_csr_address [7]),
        .O(read_data_out2_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    read_data_out2_carry_i_3
       (.I0(\processor/wb_csr_address [3]),
        .I1(\csr_addr[3]_i_1_n_0 ),
        .I2(\csr_addr[5]_i_1_n_0 ),
        .I3(\processor/wb_csr_address [5]),
        .I4(\csr_addr[4]_i_1_n_0 ),
        .I5(\processor/wb_csr_address [4]),
        .O(read_data_out2_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    read_data_out2_carry_i_4
       (.I0(\processor/wb_csr_address [0]),
        .I1(csr_addr),
        .I2(\csr_addr[2]_i_1_n_0 ),
        .I3(\processor/wb_csr_address [2]),
        .I4(\csr_addr[1]_i_1_n_0 ),
        .I5(\processor/wb_csr_address [1]),
        .O(read_data_out2_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[0]_i_1 
       (.I0(\processor/wb_csr_data [0]),
        .I1(\processor/csr_unit/read_data_out__582 [0]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(read_data_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[0]_i_2 
       (.I0(data16[0]),
        .I1(\read_data_out[0]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(read_data_out_reg),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[0]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[0]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_ ),
        .I1(data14[0]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_ ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[0]),
        .O(\read_data_out[0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \read_data_out[0]_i_5 
       (.I0(\read_data_out[31]_i_12_n_0 ),
        .I1(\read_data_out[0]_i_8_n_0 ),
        .O(\read_data_out[0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA0A0CFC0)) 
    \read_data_out[0]_i_6 
       (.I0(mbadaddr[0]),
        .I1(\processor/mie [0]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(mtvec[0]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .O(\read_data_out[0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[0]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_ ),
        .I1(mtime_compare[0]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/counter_mtime_reg [0]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data8[0]),
        .O(\read_data_out[0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[0]_i_8 
       (.I0(mepc[0]),
        .I1(mscratch[0]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/ie ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(fromhost[0]),
        .O(\read_data_out[0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[10]_i_1 
       (.I0(\processor/wb_csr_data [10]),
        .I1(\processor/csr_unit/read_data_out__582 [10]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[10]_i_2 
       (.I0(data16[10]),
        .I1(\read_data_out[10]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[10]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[10]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[10]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[10] ),
        .I1(data14[10]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[10] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[10]),
        .O(\read_data_out[10]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFCFAFC000000000)) 
    \read_data_out[10]_i_5 
       (.I0(mepc[10]),
        .I1(mscratch[10]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(fromhost[10]),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[10]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA0A0CFC0)) 
    \read_data_out[10]_i_6 
       (.I0(mbadaddr[10]),
        .I1(\processor/mie [10]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(mtvec[10]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .O(\read_data_out[10]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[10]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[10] ),
        .I1(mtime_compare[10]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [10]),
        .O(\read_data_out[10]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[11]_i_1 
       (.I0(\processor/wb_csr_data [11]),
        .I1(\processor/csr_unit/read_data_out__582 [11]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[11]_i_2 
       (.I0(data16[11]),
        .I1(\read_data_out[11]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[11]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[11]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[11]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[11] ),
        .I1(data14[11]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[11] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[11]),
        .O(\read_data_out[11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFCFAFC000000000)) 
    \read_data_out[11]_i_5 
       (.I0(mepc[11]),
        .I1(mscratch[11]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(fromhost[11]),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[11]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA0A0CFC0)) 
    \read_data_out[11]_i_6 
       (.I0(mbadaddr[11]),
        .I1(\processor/mie [11]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(mtvec[11]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .O(\read_data_out[11]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[11]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[11] ),
        .I1(mtime_compare[11]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [11]),
        .O(\read_data_out[11]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[12]_i_1 
       (.I0(\processor/wb_csr_data [12]),
        .I1(\processor/csr_unit/read_data_out__582 [12]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[12]_i_2 
       (.I0(data16[12]),
        .I1(\read_data_out[12]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[12]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[12]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[12]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[12] ),
        .I1(data14[12]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[12] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[12]),
        .O(\read_data_out[12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A0CFC000000000)) 
    \read_data_out[12]_i_5 
       (.I0(mepc[12]),
        .I1(mscratch[12]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(fromhost[12]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA0A0CFC0)) 
    \read_data_out[12]_i_6 
       (.I0(mbadaddr[12]),
        .I1(\processor/mie [12]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(mtvec[12]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .O(\read_data_out[12]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[12]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[12] ),
        .I1(mtime_compare[12]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [12]),
        .O(\read_data_out[12]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[13]_i_1 
       (.I0(\processor/wb_csr_data [13]),
        .I1(\processor/csr_unit/read_data_out__582 [13]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[13]_i_2 
       (.I0(data16[13]),
        .I1(\read_data_out[13]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[13]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[13]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[13]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[13] ),
        .I1(data14[13]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[13] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[13]),
        .O(\read_data_out[13]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A0CFC000000000)) 
    \read_data_out[13]_i_5 
       (.I0(mepc[13]),
        .I1(mscratch[13]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(fromhost[13]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[13]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA0A0CFC0)) 
    \read_data_out[13]_i_6 
       (.I0(mbadaddr[13]),
        .I1(\processor/mie [13]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(mtvec[13]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .O(\read_data_out[13]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[13]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[13] ),
        .I1(mtime_compare[13]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [13]),
        .O(\read_data_out[13]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[14]_i_1 
       (.I0(\processor/wb_csr_data [14]),
        .I1(\processor/csr_unit/read_data_out__582 [14]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[14]_i_2 
       (.I0(data16[14]),
        .I1(\read_data_out[14]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[14]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[14]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[14]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[14] ),
        .I1(data14[14]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[14] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[14]),
        .O(\read_data_out[14]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A0CFC000000000)) 
    \read_data_out[14]_i_5 
       (.I0(mepc[14]),
        .I1(mscratch[14]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(fromhost[14]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[14]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA0A0CFC0)) 
    \read_data_out[14]_i_6 
       (.I0(mbadaddr[14]),
        .I1(\processor/mie [14]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(mtvec[14]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .O(\read_data_out[14]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[14]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[14] ),
        .I1(mtime_compare[14]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [14]),
        .O(\read_data_out[14]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[15]_i_1 
       (.I0(\processor/wb_csr_data [15]),
        .I1(\processor/csr_unit/read_data_out__582 [15]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[15]_i_2 
       (.I0(data16[15]),
        .I1(\read_data_out[15]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[15]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[15]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[15]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[15] ),
        .I1(data14[15]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[15] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[15]),
        .O(\read_data_out[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF0000000CCFFAA00)) 
    \read_data_out[15]_i_5 
       (.I0(fromhost[15]),
        .I1(mscratch[15]),
        .I2(mepc[15]),
        .I3(\read_data_out[31]_i_12_n_0 ),
        .I4(\read_data_out[31]_i_8_n_0 ),
        .I5(\read_data_out[31]_i_9_n_0 ),
        .O(\read_data_out[15]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA0A0CFC0)) 
    \read_data_out[15]_i_6 
       (.I0(mbadaddr[15]),
        .I1(\processor/mie [15]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(mtvec[15]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .O(\read_data_out[15]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[15]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[15] ),
        .I1(mtime_compare[15]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [15]),
        .O(\read_data_out[15]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[16]_i_1 
       (.I0(\processor/wb_csr_data [16]),
        .I1(\processor/csr_unit/read_data_out__582 [16]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[16]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[16]_i_2 
       (.I0(data16[16]),
        .I1(\read_data_out[16]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[16]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[16]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[16]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[16] ),
        .I1(data14[16]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[16] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[16]),
        .O(\read_data_out[16]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A0CFC000000000)) 
    \read_data_out[16]_i_5 
       (.I0(mepc[16]),
        .I1(mscratch[16]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(fromhost[16]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[16]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA0A0CFC0)) 
    \read_data_out[16]_i_6 
       (.I0(mbadaddr[16]),
        .I1(\processor/mie [16]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(mtvec[16]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .O(\read_data_out[16]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[16]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[16] ),
        .I1(mtime_compare[16]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [16]),
        .O(\read_data_out[16]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[17]_i_1 
       (.I0(\processor/wb_csr_data [17]),
        .I1(\processor/csr_unit/read_data_out__582 [17]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[17]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[17]_i_2 
       (.I0(data16[17]),
        .I1(\read_data_out[17]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[17]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[17]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[17]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[17] ),
        .I1(data14[17]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[17] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[17]),
        .O(\read_data_out[17]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A0CFC000000000)) 
    \read_data_out[17]_i_5 
       (.I0(mepc[17]),
        .I1(mscratch[17]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(fromhost[17]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[17]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA0A0CFC0)) 
    \read_data_out[17]_i_6 
       (.I0(mbadaddr[17]),
        .I1(\processor/mie [17]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(mtvec[17]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .O(\read_data_out[17]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[17]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[17] ),
        .I1(mtime_compare[17]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [17]),
        .O(\read_data_out[17]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[18]_i_1 
       (.I0(\processor/wb_csr_data [18]),
        .I1(\processor/csr_unit/read_data_out__582 [18]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[18]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[18]_i_2 
       (.I0(data16[18]),
        .I1(\read_data_out[18]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[18]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[18]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[18]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[18] ),
        .I1(data14[18]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[18] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[18]),
        .O(\read_data_out[18]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A0CFC000000000)) 
    \read_data_out[18]_i_5 
       (.I0(mepc[18]),
        .I1(mscratch[18]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(fromhost[18]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[18]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA0A0CFC0)) 
    \read_data_out[18]_i_6 
       (.I0(mbadaddr[18]),
        .I1(\processor/mie [18]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(mtvec[18]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .O(\read_data_out[18]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[18]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[18] ),
        .I1(mtime_compare[18]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [18]),
        .O(\read_data_out[18]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[19]_i_1 
       (.I0(\processor/wb_csr_data [19]),
        .I1(\processor/csr_unit/read_data_out__582 [19]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[19]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[19]_i_2 
       (.I0(data16[19]),
        .I1(\read_data_out[19]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[19]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[19]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[19]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[19] ),
        .I1(data14[19]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[19] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[19]),
        .O(\read_data_out[19]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A0CFC000000000)) 
    \read_data_out[19]_i_5 
       (.I0(mepc[19]),
        .I1(mscratch[19]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(fromhost[19]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[19]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA0A0CFC0)) 
    \read_data_out[19]_i_6 
       (.I0(mbadaddr[19]),
        .I1(\processor/mie [19]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(mtvec[19]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .O(\read_data_out[19]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[19]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[19] ),
        .I1(mtime_compare[19]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [19]),
        .O(\read_data_out[19]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[1]_i_1 
       (.I0(\processor/wb_csr_data [1]),
        .I1(\processor/csr_unit/read_data_out__582 [1]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[1]_i_2 
       (.I0(data16[1]),
        .I1(\read_data_out[1]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[1]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[1]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[1]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[1] ),
        .I1(data14[1]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[1] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[1]),
        .O(\read_data_out[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFCFAFC000000000)) 
    \read_data_out[1]_i_5 
       (.I0(mepc[1]),
        .I1(mscratch[1]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(fromhost[1]),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA0A0CFC0)) 
    \read_data_out[1]_i_6 
       (.I0(mbadaddr[1]),
        .I1(\processor/mie [1]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(mtvec[1]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .O(\read_data_out[1]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[1]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[1] ),
        .I1(mtime_compare[1]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/counter_mtime_reg [1]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data8[1]),
        .O(\read_data_out[1]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[20]_i_1 
       (.I0(\processor/wb_csr_data [20]),
        .I1(\processor/csr_unit/read_data_out__582 [20]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[20]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[20]_i_2 
       (.I0(data16[20]),
        .I1(\read_data_out[20]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[20]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[20]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[20]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[20] ),
        .I1(data14[20]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[20] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[20]),
        .O(\read_data_out[20]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A0CFC000000000)) 
    \read_data_out[20]_i_5 
       (.I0(mepc[20]),
        .I1(mscratch[20]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(fromhost[20]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[20]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA0A0CFC0)) 
    \read_data_out[20]_i_6 
       (.I0(mbadaddr[20]),
        .I1(\processor/mie [20]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(mtvec[20]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .O(\read_data_out[20]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[20]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[20] ),
        .I1(mtime_compare[20]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [20]),
        .O(\read_data_out[20]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[21]_i_1 
       (.I0(\processor/wb_csr_data [21]),
        .I1(\processor/csr_unit/read_data_out__582 [21]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[21]_i_2 
       (.I0(data16[21]),
        .I1(\read_data_out[21]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[21]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[21]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[21]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[21] ),
        .I1(data14[21]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[21] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[21]),
        .O(\read_data_out[21]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A0CFC000000000)) 
    \read_data_out[21]_i_5 
       (.I0(mepc[21]),
        .I1(mscratch[21]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(fromhost[21]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[21]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA0A0CFC0)) 
    \read_data_out[21]_i_6 
       (.I0(mbadaddr[21]),
        .I1(\processor/mie [21]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(mtvec[21]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .O(\read_data_out[21]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[21]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[21] ),
        .I1(mtime_compare[21]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [21]),
        .O(\read_data_out[21]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[22]_i_1 
       (.I0(\processor/wb_csr_data [22]),
        .I1(\processor/csr_unit/read_data_out__582 [22]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[22]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[22]_i_2 
       (.I0(data16[22]),
        .I1(\read_data_out[22]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[22]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[22]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[22]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[22] ),
        .I1(data14[22]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[22] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[22]),
        .O(\read_data_out[22]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A0CFC000000000)) 
    \read_data_out[22]_i_5 
       (.I0(mepc[22]),
        .I1(mscratch[22]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(fromhost[22]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[22]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA0A0CFC0)) 
    \read_data_out[22]_i_6 
       (.I0(mbadaddr[22]),
        .I1(\processor/mie [22]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(mtvec[22]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .O(\read_data_out[22]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[22]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[22] ),
        .I1(mtime_compare[22]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [22]),
        .O(\read_data_out[22]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[23]_i_1 
       (.I0(\processor/wb_csr_data [23]),
        .I1(\processor/csr_unit/read_data_out__582 [23]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[23]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[23]_i_2 
       (.I0(data16[23]),
        .I1(\read_data_out[23]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[23]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[23]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[23]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[23] ),
        .I1(data14[23]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[23] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[23]),
        .O(\read_data_out[23]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A0CFC000000000)) 
    \read_data_out[23]_i_5 
       (.I0(mepc[23]),
        .I1(mscratch[23]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(fromhost[23]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[23]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA0A0CFC0)) 
    \read_data_out[23]_i_6 
       (.I0(mbadaddr[23]),
        .I1(\processor/mie [23]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(mtvec[23]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .O(\read_data_out[23]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[23]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[23] ),
        .I1(mtime_compare[23]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [23]),
        .O(\read_data_out[23]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[24]_i_1 
       (.I0(\processor/wb_csr_data [24]),
        .I1(\processor/csr_unit/read_data_out__582 [24]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[24]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[24]_i_2 
       (.I0(data16[24]),
        .I1(\read_data_out[24]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[24]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[24]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[24]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[24] ),
        .I1(data14[24]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[24] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[24]),
        .O(\read_data_out[24]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A0CFC000000000)) 
    \read_data_out[24]_i_5 
       (.I0(mepc[24]),
        .I1(mscratch[24]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(fromhost[24]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[24]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[24]_i_6 
       (.I0(mbadaddr[24]),
        .I1(\processor/mie [24]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(irq[0]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(mtvec[24]),
        .O(\read_data_out[24]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[24]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[24] ),
        .I1(mtime_compare[24]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [24]),
        .O(\read_data_out[24]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[25]_i_1 
       (.I0(\processor/wb_csr_data [25]),
        .I1(\processor/csr_unit/read_data_out__582 [25]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[25]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[25]_i_2 
       (.I0(data16[25]),
        .I1(\read_data_out[25]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[25]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[25]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[25]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[25] ),
        .I1(data14[25]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[25] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[25]),
        .O(\read_data_out[25]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A0CFC000000000)) 
    \read_data_out[25]_i_5 
       (.I0(mepc[25]),
        .I1(mscratch[25]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(fromhost[25]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[25]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[25]_i_6 
       (.I0(mbadaddr[25]),
        .I1(\processor/mie [25]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(irq[1]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(mtvec[25]),
        .O(\read_data_out[25]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[25]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[25] ),
        .I1(mtime_compare[25]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [25]),
        .O(\read_data_out[25]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[26]_i_1 
       (.I0(\processor/wb_csr_data [26]),
        .I1(\processor/csr_unit/read_data_out__582 [26]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[26]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[26]_i_2 
       (.I0(data16[26]),
        .I1(\read_data_out[26]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[26]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[26]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[26]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[26] ),
        .I1(data14[26]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[26] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[26]),
        .O(\read_data_out[26]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A0CFC000000000)) 
    \read_data_out[26]_i_5 
       (.I0(mepc[26]),
        .I1(mscratch[26]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(fromhost[26]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[26]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[26]_i_6 
       (.I0(mbadaddr[26]),
        .I1(\processor/mie [26]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(irq[2]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(mtvec[26]),
        .O(\read_data_out[26]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[26]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[26] ),
        .I1(mtime_compare[26]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [26]),
        .O(\read_data_out[26]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[27]_i_1 
       (.I0(\processor/wb_csr_data [27]),
        .I1(\processor/csr_unit/read_data_out__582 [27]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[27]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[27]_i_2 
       (.I0(data16[27]),
        .I1(\read_data_out[27]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[27]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[27]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[27]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[27] ),
        .I1(data14[27]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[27] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[27]),
        .O(\read_data_out[27]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A0CFC000000000)) 
    \read_data_out[27]_i_5 
       (.I0(mepc[27]),
        .I1(mscratch[27]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(fromhost[27]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[27]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[27]_i_6 
       (.I0(mbadaddr[27]),
        .I1(\processor/mie [27]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(irq[3]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(mtvec[27]),
        .O(\read_data_out[27]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[27]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[27] ),
        .I1(mtime_compare[27]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [27]),
        .O(\read_data_out[27]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[28]_i_1 
       (.I0(\processor/wb_csr_data [28]),
        .I1(\processor/csr_unit/read_data_out__582 [28]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[28]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[28]_i_2 
       (.I0(data16[28]),
        .I1(\read_data_out[28]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[28]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[28]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[28]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[28] ),
        .I1(data14[28]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[28] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[28]),
        .O(\read_data_out[28]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A0CFC000000000)) 
    \read_data_out[28]_i_5 
       (.I0(mepc[28]),
        .I1(mscratch[28]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(fromhost[28]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[28]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[28]_i_6 
       (.I0(mbadaddr[28]),
        .I1(\processor/mie [28]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(irq[4]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(mtvec[28]),
        .O(\read_data_out[28]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[28]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[28] ),
        .I1(mtime_compare[28]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [28]),
        .O(\read_data_out[28]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[29]_i_1 
       (.I0(\processor/wb_csr_data [29]),
        .I1(\processor/csr_unit/read_data_out__582 [29]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[29]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[29]_i_2 
       (.I0(data16[29]),
        .I1(\read_data_out[29]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[29]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[29]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[29]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[29] ),
        .I1(data14[29]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[29] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[29]),
        .O(\read_data_out[29]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A0CFC000000000)) 
    \read_data_out[29]_i_5 
       (.I0(mepc[29]),
        .I1(mscratch[29]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(fromhost[29]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[29]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[29]_i_6 
       (.I0(mbadaddr[29]),
        .I1(\processor/mie [29]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(irq[5]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(mtvec[29]),
        .O(\read_data_out[29]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[29]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[29] ),
        .I1(mtime_compare[29]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [29]),
        .O(\read_data_out[29]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[2]_i_1 
       (.I0(\processor/wb_csr_data [2]),
        .I1(\processor/csr_unit/read_data_out__582 [2]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[2]_i_2 
       (.I0(data16[2]),
        .I1(\read_data_out[2]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[2]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[2]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[2]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[2] ),
        .I1(data14[2]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[2] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[2]),
        .O(\read_data_out[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFCFAFC000000000)) 
    \read_data_out[2]_i_5 
       (.I0(mepc[2]),
        .I1(mscratch[2]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(fromhost[2]),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA0A0CFC0)) 
    \read_data_out[2]_i_6 
       (.I0(mbadaddr[2]),
        .I1(\processor/mie [2]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(mtvec[2]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .O(\read_data_out[2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[2]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[2] ),
        .I1(mtime_compare[2]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/counter_mtime_reg [2]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data8[2]),
        .O(\read_data_out[2]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[30]_i_1 
       (.I0(\processor/wb_csr_data [30]),
        .I1(\processor/csr_unit/read_data_out__582 [30]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[30]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[30]_i_2 
       (.I0(data16[30]),
        .I1(\read_data_out[30]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[30]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[30]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[30]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[30] ),
        .I1(data14[30]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[30] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[30]),
        .O(\read_data_out[30]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A0CFC000000000)) 
    \read_data_out[30]_i_5 
       (.I0(mepc[30]),
        .I1(mscratch[30]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(fromhost[30]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[30]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[30]_i_6 
       (.I0(mbadaddr[30]),
        .I1(\processor/mie [30]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(irq[6]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(mtvec[30]),
        .O(\read_data_out[30]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[30]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[30] ),
        .I1(mtime_compare[30]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [30]),
        .O(\read_data_out[30]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[31]_i_1 
       (.I0(\processor/wb_csr_data [31]),
        .I1(\processor/csr_unit/read_data_out__582 [31]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \read_data_out[31]_i_10 
       (.I0(\csr_addr[2]_i_1_n_0 ),
        .I1(\csr_addr[3]_i_1_n_0 ),
        .O(\read_data_out[31]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFDFFFDFDFDFFFDF)) 
    \read_data_out[31]_i_11 
       (.I0(\csr_addr[11]_i_1_n_0 ),
        .I1(\csr_addr[4]_i_1_n_0 ),
        .I2(\csr_addr[10]_i_1_n_0 ),
        .I3(csr_addr),
        .I4(\csr_addr[7]_i_1_n_0 ),
        .I5(\csr_addr[1]_i_1_n_0 ),
        .O(\read_data_out[31]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000200020002AA02)) 
    \read_data_out[31]_i_12 
       (.I0(\read_data_out[31]_i_20_n_0 ),
        .I1(\read_data_out[31]_i_21_n_0 ),
        .I2(\csr_addr[5]_i_1_n_0 ),
        .I3(csr_addr),
        .I4(\read_data_out[31]_i_22_n_0 ),
        .I5(\csr_addr[1]_i_1_n_0 ),
        .O(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[31]_i_13 
       (.I0(mbadaddr[31]),
        .I1(\processor/mie [31]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(irq[7]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(mtvec[31]),
        .O(\read_data_out[31]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[31]_i_14 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[31] ),
        .I1(mtime_compare[31]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/counter_mtime_reg [31]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data8[31]),
        .O(\read_data_out[31]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000110)) 
    \read_data_out[31]_i_15 
       (.I0(\csr_addr[3]_i_1_n_0 ),
        .I1(\csr_addr[7]_i_1_n_0 ),
        .I2(\csr_addr[9]_i_1_n_0 ),
        .I3(\csr_addr[11]_i_1_n_0 ),
        .I4(\csr_addr[4]_i_1_n_0 ),
        .O(\read_data_out[31]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1070000400000000)) 
    \read_data_out[31]_i_16 
       (.I0(\csr_addr[6]_i_1_n_0 ),
        .I1(\csr_addr[10]_i_1_n_0 ),
        .I2(\csr_addr[9]_i_1_n_0 ),
        .I3(\csr_addr[5]_i_1_n_0 ),
        .I4(\csr_addr[8]_i_1_n_0 ),
        .I5(\read_data_out[31]_i_23_n_0 ),
        .O(\read_data_out[31]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFC6)) 
    \read_data_out[31]_i_17 
       (.I0(\csr_addr[6]_i_1_n_0 ),
        .I1(\csr_addr[2]_i_1_n_0 ),
        .I2(\csr_addr[1]_i_1_n_0 ),
        .I3(\read_data_out[31]_i_24_n_0 ),
        .I4(\csr_addr[4]_i_1_n_0 ),
        .I5(\csr_addr[3]_i_1_n_0 ),
        .O(\read_data_out[31]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFA656)) 
    \read_data_out[31]_i_18 
       (.I0(\csr_addr[11]_i_1_n_0 ),
        .I1(\csr_addr[10]_i_1_n_0 ),
        .I2(csr_addr),
        .I3(\csr_addr[8]_i_1_n_0 ),
        .I4(\read_data_out[31]_i_25_n_0 ),
        .O(\read_data_out[31]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEE1011)) 
    \read_data_out[31]_i_19 
       (.I0(\csr_addr[6]_i_1_n_0 ),
        .I1(\csr_addr[2]_i_1_n_0 ),
        .I2(\csr_addr[8]_i_1_n_0 ),
        .I3(\csr_addr[7]_i_1_n_0 ),
        .I4(csr_addr),
        .I5(\read_data_out[31]_i_26_n_0 ),
        .O(\read_data_out[31]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[31]_i_2 
       (.I0(data16[31]),
        .I1(\read_data_out[31]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[31]_i_5_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[31]_i_7_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000110)) 
    \read_data_out[31]_i_20 
       (.I0(\csr_addr[2]_i_1_n_0 ),
        .I1(\csr_addr[4]_i_1_n_0 ),
        .I2(\csr_addr[9]_i_1_n_0 ),
        .I3(\csr_addr[11]_i_1_n_0 ),
        .I4(\csr_addr[3]_i_1_n_0 ),
        .O(\read_data_out[31]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFDFFFFBFFDFFFDFF)) 
    \read_data_out[31]_i_21 
       (.I0(\csr_addr[9]_i_1_n_0 ),
        .I1(\csr_addr[10]_i_1_n_0 ),
        .I2(\csr_addr[7]_i_1_n_0 ),
        .I3(\csr_addr[8]_i_1_n_0 ),
        .I4(\csr_addr[6]_i_1_n_0 ),
        .I5(\csr_addr[1]_i_1_n_0 ),
        .O(\read_data_out[31]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFBFFBB7FFFFFFEF)) 
    \read_data_out[31]_i_22 
       (.I0(\csr_addr[5]_i_1_n_0 ),
        .I1(\csr_addr[9]_i_1_n_0 ),
        .I2(\csr_addr[10]_i_1_n_0 ),
        .I3(\csr_addr[6]_i_1_n_0 ),
        .I4(\csr_addr[7]_i_1_n_0 ),
        .I5(\csr_addr[8]_i_1_n_0 ),
        .O(\read_data_out[31]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0050005000980598)) 
    \read_data_out[31]_i_23 
       (.I0(\csr_addr[1]_i_1_n_0 ),
        .I1(\csr_addr[6]_i_1_n_0 ),
        .I2(csr_addr),
        .I3(\csr_addr[2]_i_1_n_0 ),
        .I4(\csr_addr[10]_i_1_n_0 ),
        .I5(\csr_addr[5]_i_1_n_0 ),
        .O(\read_data_out[31]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFCFFFFFD)) 
    \read_data_out[31]_i_24 
       (.I0(\csr_addr[10]_i_1_n_0 ),
        .I1(\csr_addr[5]_i_1_n_0 ),
        .I2(\read_data_out[31]_i_27_n_0 ),
        .I3(\csr_addr[8]_i_1_n_0 ),
        .I4(\csr_addr[9]_i_1_n_0 ),
        .O(\read_data_out[31]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00FF00FDFFFD00)) 
    \read_data_out[31]_i_25 
       (.I0(\csr_addr[8]_i_1_n_0 ),
        .I1(\csr_addr[10]_i_1_n_0 ),
        .I2(csr_addr),
        .I3(\csr_addr[6]_i_1_n_0 ),
        .I4(\csr_addr[1]_i_1_n_0 ),
        .I5(\csr_addr[7]_i_1_n_0 ),
        .O(\read_data_out[31]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFBF00000000)) 
    \read_data_out[31]_i_26 
       (.I0(\read_data_out[31]_i_28_n_0 ),
        .I1(\csr_addr[8]_i_1_n_0 ),
        .I2(\csr_addr[9]_i_1_n_0 ),
        .I3(\csr_addr[11]_i_1_n_0 ),
        .I4(\csr_addr[10]_i_1_n_0 ),
        .I5(\read_data_out[31]_i_29_n_0 ),
        .O(\read_data_out[31]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h82)) 
    \read_data_out[31]_i_27 
       (.I0(\csr_addr[7]_i_1_n_0 ),
        .I1(\csr_addr[1]_i_1_n_0 ),
        .I2(csr_addr),
        .O(\read_data_out[31]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \read_data_out[31]_i_28 
       (.I0(\csr_addr[4]_i_1_n_0 ),
        .I1(\csr_addr[7]_i_1_n_0 ),
        .I2(\csr_addr[2]_i_1_n_0 ),
        .I3(\csr_addr[3]_i_1_n_0 ),
        .O(\read_data_out[31]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAA22AAAAA8AAA)) 
    \read_data_out[31]_i_29 
       (.I0(\read_data_out[31]_i_30_n_0 ),
        .I1(\csr_addr[8]_i_1_n_0 ),
        .I2(\csr_addr[11]_i_1_n_0 ),
        .I3(\csr_addr[7]_i_1_n_0 ),
        .I4(\read_data_out[31]_i_31_n_0 ),
        .I5(\csr_addr[9]_i_1_n_0 ),
        .O(\read_data_out[31]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[31]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[31] ),
        .I1(data14[31]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[31] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[31]),
        .O(\read_data_out[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    \read_data_out[31]_i_30 
       (.I0(\read_data_out[31]_i_32_n_0 ),
        .I1(\csr_addr[6]_i_1_n_0 ),
        .I2(\read_data_out[31]_i_33_n_0 ),
        .I3(\csr_addr[7]_i_1_n_0 ),
        .I4(\csr_addr[11]_i_1_n_0 ),
        .I5(\csr_addr[9]_i_1_n_0 ),
        .O(\read_data_out[31]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFD)) 
    \read_data_out[31]_i_31 
       (.I0(\csr_addr[10]_i_1_n_0 ),
        .I1(\csr_addr[3]_i_1_n_0 ),
        .I2(\csr_addr[2]_i_1_n_0 ),
        .I3(\csr_addr[6]_i_1_n_0 ),
        .I4(\csr_addr[4]_i_1_n_0 ),
        .O(\read_data_out[31]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \read_data_out[31]_i_32 
       (.I0(\csr_addr[4]_i_1_n_0 ),
        .I1(\csr_addr[3]_i_1_n_0 ),
        .O(\read_data_out[31]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \read_data_out[31]_i_33 
       (.I0(\csr_addr[10]_i_1_n_0 ),
        .I1(\csr_addr[8]_i_1_n_0 ),
        .O(\read_data_out[31]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \read_data_out[31]_i_4 
       (.I0(\read_data_out[31]_i_10_n_0 ),
        .I1(\read_data_out[31]_i_11_n_0 ),
        .I2(\csr_addr[8]_i_1_n_0 ),
        .I3(\csr_addr[9]_i_1_n_0 ),
        .I4(\csr_addr[5]_i_1_n_0 ),
        .I5(\csr_addr[6]_i_1_n_0 ),
        .O(\read_data_out[31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB888)) 
    \read_data_out[31]_i_6 
       (.I0(\read_data_out[31]_i_12_n_0 ),
        .I1(\read_data_out[31]_i_4_n_0 ),
        .I2(\read_data_out[31]_i_15_n_0 ),
        .I3(\read_data_out[31]_i_16_n_0 ),
        .O(\read_data_out[31]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A0CFC000000000)) 
    \read_data_out[31]_i_7 
       (.I0(mepc[31]),
        .I1(mscratch[31]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(fromhost[31]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[31]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4C31)) 
    \read_data_out[31]_i_8 
       (.I0(\csr_addr[10]_i_1_n_0 ),
        .I1(\csr_addr[7]_i_1_n_0 ),
        .I2(csr_addr),
        .I3(\csr_addr[8]_i_1_n_0 ),
        .I4(\read_data_out[31]_i_17_n_0 ),
        .I5(\read_data_out[31]_i_18_n_0 ),
        .O(\read_data_out[31]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA8AFA8)) 
    \read_data_out[31]_i_9 
       (.I0(\csr_addr[1]_i_1_n_0 ),
        .I1(\csr_addr[2]_i_1_n_0 ),
        .I2(csr_addr),
        .I3(\csr_addr[5]_i_1_n_0 ),
        .I4(\csr_addr[10]_i_1_n_0 ),
        .I5(\read_data_out[31]_i_19_n_0 ),
        .O(\read_data_out[31]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[3]_i_1 
       (.I0(\processor/wb_csr_data [3]),
        .I1(\processor/csr_unit/read_data_out__582 [3]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[3]_i_2 
       (.I0(data16[3]),
        .I1(\read_data_out[3]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[3]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[3]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[3]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[3] ),
        .I1(data14[3]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[3] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[3]),
        .O(\read_data_out[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \read_data_out[3]_i_5 
       (.I0(\read_data_out[31]_i_12_n_0 ),
        .I1(\read_data_out[3]_i_8_n_0 ),
        .O(\read_data_out[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[3]_i_6 
       (.I0(mbadaddr[3]),
        .I1(\processor/mie [3]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/software_interrupt ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(mtvec[3]),
        .O(\read_data_out[3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[3]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[3] ),
        .I1(mtime_compare[3]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/counter_mtime_reg [3]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data8[3]),
        .O(\read_data_out[3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[3]_i_8 
       (.I0(mepc[3]),
        .I1(mscratch[3]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/ie1 ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(fromhost[3]),
        .O(\read_data_out[3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[4]_i_1 
       (.I0(\processor/wb_csr_data [4]),
        .I1(\processor/csr_unit/read_data_out__582 [4]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[4]_i_2 
       (.I0(data16[4]),
        .I1(\read_data_out[4]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[4]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[4]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[4]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[4] ),
        .I1(data14[4]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[4] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[4]),
        .O(\read_data_out[4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFCFAFC000000000)) 
    \read_data_out[4]_i_5 
       (.I0(mepc[4]),
        .I1(mscratch[4]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(fromhost[4]),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA0A0CFC0)) 
    \read_data_out[4]_i_6 
       (.I0(mbadaddr[4]),
        .I1(\processor/mie [4]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(mtvec[4]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .O(\read_data_out[4]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[4]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[4] ),
        .I1(mtime_compare[4]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/counter_mtime_reg [4]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data8[4]),
        .O(\read_data_out[4]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[5]_i_1 
       (.I0(\processor/wb_csr_data [5]),
        .I1(\processor/csr_unit/read_data_out__582 [5]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[5]_i_2 
       (.I0(data16[5]),
        .I1(\read_data_out[5]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[5]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[5]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[5]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[5] ),
        .I1(data14[5]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[5] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[5]),
        .O(\read_data_out[5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFCFAFC000000000)) 
    \read_data_out[5]_i_5 
       (.I0(mepc[5]),
        .I1(mscratch[5]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(fromhost[5]),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[5]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA0A0CFC0)) 
    \read_data_out[5]_i_6 
       (.I0(mbadaddr[5]),
        .I1(\processor/mie [5]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(mtvec[5]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .O(\read_data_out[5]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[5]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[5] ),
        .I1(mtime_compare[5]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [5]),
        .O(\read_data_out[5]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[6]_i_1 
       (.I0(\processor/wb_csr_data [6]),
        .I1(\processor/csr_unit/read_data_out__582 [6]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[6]_i_2 
       (.I0(data16[6]),
        .I1(\read_data_out[6]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[6]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[6]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[6]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[6] ),
        .I1(data14[6]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[6] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[6]),
        .O(\read_data_out[6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A0CFC000000000)) 
    \read_data_out[6]_i_5 
       (.I0(mepc[6]),
        .I1(mscratch[6]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(fromhost[6]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[6]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA0A0CFC0)) 
    \read_data_out[6]_i_6 
       (.I0(mbadaddr[6]),
        .I1(\processor/mie [6]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(mtvec[6]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .O(\read_data_out[6]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[6]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[6] ),
        .I1(mtime_compare[6]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [6]),
        .O(\read_data_out[6]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[7]_i_1 
       (.I0(\processor/wb_csr_data [7]),
        .I1(\processor/csr_unit/read_data_out__582 [7]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[7]_i_2 
       (.I0(data16[7]),
        .I1(\read_data_out[7]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[7]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[7]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[7]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[7] ),
        .I1(data14[7]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[7] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[7]),
        .O(\read_data_out[7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFCFAFC000000000)) 
    \read_data_out[7]_i_5 
       (.I0(mepc[7]),
        .I1(mscratch[7]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(fromhost[7]),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[7]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[7]_i_6 
       (.I0(mbadaddr[7]),
        .I1(\processor/mie [7]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/timer_interrupt ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(mtvec[7]),
        .O(\read_data_out[7]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[7]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[7] ),
        .I1(mtime_compare[7]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [7]),
        .O(\read_data_out[7]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[8]_i_1 
       (.I0(\processor/wb_csr_data [8]),
        .I1(\processor/csr_unit/read_data_out__582 [8]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[8]_i_2 
       (.I0(data16[8]),
        .I1(\read_data_out[8]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[8]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[8]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[8]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[8] ),
        .I1(data14[8]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[8] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[8]),
        .O(\read_data_out[8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBB3BB333B939B131)) 
    \read_data_out[8]_i_5 
       (.I0(\read_data_out[31]_i_12_n_0 ),
        .I1(\read_data_out[31]_i_8_n_0 ),
        .I2(\read_data_out[31]_i_9_n_0 ),
        .I3(mepc[8]),
        .I4(mscratch[8]),
        .I5(fromhost[8]),
        .O(\read_data_out[8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA0A0CFC0)) 
    \read_data_out[8]_i_6 
       (.I0(mbadaddr[8]),
        .I1(\processor/mie [8]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(mtvec[8]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .O(\read_data_out[8]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[8]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[8] ),
        .I1(mtime_compare[8]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [8]),
        .O(\read_data_out[8]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAACCCCC)) 
    \read_data_out[9]_i_1 
       (.I0(\processor/wb_csr_data [9]),
        .I1(\processor/csr_unit/read_data_out__582 [9]),
        .I2(\processor/wb_csr_write [0]),
        .I3(\processor/wb_csr_write [1]),
        .I4(\processor/csr_unit/read_data_out2__3 ),
        .O(\read_data_out[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[9]_i_2 
       (.I0(data16[9]),
        .I1(\read_data_out[9]_i_3_n_0 ),
        .I2(\read_data_out[31]_i_4_n_0 ),
        .I3(\read_data_out_reg[9]_i_4_n_0 ),
        .I4(\read_data_out[31]_i_6_n_0 ),
        .I5(\read_data_out[9]_i_5_n_0 ),
        .O(\processor/csr_unit/read_data_out__582 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \read_data_out[9]_i_3 
       (.I0(\processor/csr_unit/instret_counter/current_count_reg_n_0_[9] ),
        .I1(data14[9]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\processor/csr_unit/cycle_counter/current_count_reg_n_0_[9] ),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(data12[9]),
        .O(\read_data_out[9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A0CFC000000000)) 
    \read_data_out[9]_i_5 
       (.I0(mepc[9]),
        .I1(mscratch[9]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(fromhost[9]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .I5(\read_data_out[31]_i_12_n_0 ),
        .O(\read_data_out[9]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA0A0CFC0)) 
    \read_data_out[9]_i_6 
       (.I0(mbadaddr[9]),
        .I1(\processor/mie [9]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(mtvec[9]),
        .I4(\read_data_out[31]_i_9_n_0 ),
        .O(\read_data_out[9]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \read_data_out[9]_i_7 
       (.I0(\processor/csr_unit/timer_counter/current_count_reg_n_0_[9] ),
        .I1(mtime_compare[9]),
        .I2(\read_data_out[31]_i_8_n_0 ),
        .I3(\read_data_out[31]_i_9_n_0 ),
        .I4(\processor/csr_unit/counter_mtime_reg [9]),
        .O(\read_data_out[9]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[0]_i_4 
       (.I0(\read_data_out[0]_i_6_n_0 ),
        .I1(\read_data_out[0]_i_7_n_0 ),
        .O(read_data_out_reg),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[10]_i_4 
       (.I0(\read_data_out[10]_i_6_n_0 ),
        .I1(\read_data_out[10]_i_7_n_0 ),
        .O(\read_data_out_reg[10]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[11]_i_4 
       (.I0(\read_data_out[11]_i_6_n_0 ),
        .I1(\read_data_out[11]_i_7_n_0 ),
        .O(\read_data_out_reg[11]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[12]_i_4 
       (.I0(\read_data_out[12]_i_6_n_0 ),
        .I1(\read_data_out[12]_i_7_n_0 ),
        .O(\read_data_out_reg[12]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[13]_i_4 
       (.I0(\read_data_out[13]_i_6_n_0 ),
        .I1(\read_data_out[13]_i_7_n_0 ),
        .O(\read_data_out_reg[13]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[14]_i_4 
       (.I0(\read_data_out[14]_i_6_n_0 ),
        .I1(\read_data_out[14]_i_7_n_0 ),
        .O(\read_data_out_reg[14]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[15]_i_4 
       (.I0(\read_data_out[15]_i_6_n_0 ),
        .I1(\read_data_out[15]_i_7_n_0 ),
        .O(\read_data_out_reg[15]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[16]_i_4 
       (.I0(\read_data_out[16]_i_6_n_0 ),
        .I1(\read_data_out[16]_i_7_n_0 ),
        .O(\read_data_out_reg[16]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[17]_i_4 
       (.I0(\read_data_out[17]_i_6_n_0 ),
        .I1(\read_data_out[17]_i_7_n_0 ),
        .O(\read_data_out_reg[17]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[18]_i_4 
       (.I0(\read_data_out[18]_i_6_n_0 ),
        .I1(\read_data_out[18]_i_7_n_0 ),
        .O(\read_data_out_reg[18]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[19]_i_4 
       (.I0(\read_data_out[19]_i_6_n_0 ),
        .I1(\read_data_out[19]_i_7_n_0 ),
        .O(\read_data_out_reg[19]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[1]_i_4 
       (.I0(\read_data_out[1]_i_6_n_0 ),
        .I1(\read_data_out[1]_i_7_n_0 ),
        .O(\read_data_out_reg[1]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[20]_i_4 
       (.I0(\read_data_out[20]_i_6_n_0 ),
        .I1(\read_data_out[20]_i_7_n_0 ),
        .O(\read_data_out_reg[20]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[21]_i_4 
       (.I0(\read_data_out[21]_i_6_n_0 ),
        .I1(\read_data_out[21]_i_7_n_0 ),
        .O(\read_data_out_reg[21]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[22]_i_4 
       (.I0(\read_data_out[22]_i_6_n_0 ),
        .I1(\read_data_out[22]_i_7_n_0 ),
        .O(\read_data_out_reg[22]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[23]_i_4 
       (.I0(\read_data_out[23]_i_6_n_0 ),
        .I1(\read_data_out[23]_i_7_n_0 ),
        .O(\read_data_out_reg[23]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[24]_i_4 
       (.I0(\read_data_out[24]_i_6_n_0 ),
        .I1(\read_data_out[24]_i_7_n_0 ),
        .O(\read_data_out_reg[24]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[25]_i_4 
       (.I0(\read_data_out[25]_i_6_n_0 ),
        .I1(\read_data_out[25]_i_7_n_0 ),
        .O(\read_data_out_reg[25]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[26]_i_4 
       (.I0(\read_data_out[26]_i_6_n_0 ),
        .I1(\read_data_out[26]_i_7_n_0 ),
        .O(\read_data_out_reg[26]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[27]_i_4 
       (.I0(\read_data_out[27]_i_6_n_0 ),
        .I1(\read_data_out[27]_i_7_n_0 ),
        .O(\read_data_out_reg[27]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[28]_i_4 
       (.I0(\read_data_out[28]_i_6_n_0 ),
        .I1(\read_data_out[28]_i_7_n_0 ),
        .O(\read_data_out_reg[28]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[29]_i_4 
       (.I0(\read_data_out[29]_i_6_n_0 ),
        .I1(\read_data_out[29]_i_7_n_0 ),
        .O(\read_data_out_reg[29]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[2]_i_4 
       (.I0(\read_data_out[2]_i_6_n_0 ),
        .I1(\read_data_out[2]_i_7_n_0 ),
        .O(\read_data_out_reg[2]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[30]_i_4 
       (.I0(\read_data_out[30]_i_6_n_0 ),
        .I1(\read_data_out[30]_i_7_n_0 ),
        .O(\read_data_out_reg[30]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[31]_i_5 
       (.I0(\read_data_out[31]_i_13_n_0 ),
        .I1(\read_data_out[31]_i_14_n_0 ),
        .O(\read_data_out_reg[31]_i_5_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[3]_i_4 
       (.I0(\read_data_out[3]_i_6_n_0 ),
        .I1(\read_data_out[3]_i_7_n_0 ),
        .O(\read_data_out_reg[3]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[4]_i_4 
       (.I0(\read_data_out[4]_i_6_n_0 ),
        .I1(\read_data_out[4]_i_7_n_0 ),
        .O(\read_data_out_reg[4]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[5]_i_4 
       (.I0(\read_data_out[5]_i_6_n_0 ),
        .I1(\read_data_out[5]_i_7_n_0 ),
        .O(\read_data_out_reg[5]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[6]_i_4 
       (.I0(\read_data_out[6]_i_6_n_0 ),
        .I1(\read_data_out[6]_i_7_n_0 ),
        .O(\read_data_out_reg[6]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[7]_i_4 
       (.I0(\read_data_out[7]_i_6_n_0 ),
        .I1(\read_data_out[7]_i_7_n_0 ),
        .O(\read_data_out_reg[7]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[8]_i_4 
       (.I0(\read_data_out[8]_i_6_n_0 ),
        .I1(\read_data_out[8]_i_7_n_0 ),
        .O(\read_data_out_reg[8]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \read_data_out_reg[9]_i_4 
       (.I0(\read_data_out[9]_i_6_n_0 ),
        .I1(\read_data_out[9]_i_7_n_0 ),
        .O(\read_data_out_reg[9]_i_4_n_0 ),
        .S(\read_data_out[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAA8)) 
    registers_reg_r1_0_31_0_5_i_1
       (.I0(\processor/wb_rd_write ),
        .I1(\processor/wb_rd_address [4]),
        .I2(\processor/wb_rd_address [3]),
        .I3(\processor/wb_rd_address [1]),
        .I4(\processor/wb_rd_address [0]),
        .I5(\processor/wb_rd_address [2]),
        .O(\processor/regfile/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h41000041)) 
    registers_reg_r1_0_31_0_5_i_10
       (.I0(registers_reg_r1_0_31_0_5_i_14_n_0),
        .I1(\processor/mem_rd_address [4]),
        .I2(\processor/execute/rs1_addr [4]),
        .I3(\processor/execute/rs1_addr [3]),
        .I4(\processor/mem_rd_address [3]),
        .O(registers_reg_r1_0_31_0_5_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    registers_reg_r1_0_31_0_5_i_11
       (.I0(\processor/execute/rs1_addr [3]),
        .I1(\processor/execute/rs1_addr [0]),
        .I2(\processor/execute/rs1_addr [2]),
        .I3(\processor/execute/rs1_addr [4]),
        .I4(\processor/execute/rs1_addr [1]),
        .O(registers_reg_r1_0_31_0_5_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h09000009)) 
    registers_reg_r1_0_31_0_5_i_12
       (.I0(\processor/execute/rs2_addr [3]),
        .I1(\processor/mem_rd_address [3]),
        .I2(\dmem_data_out_p[31]_i_5_n_0 ),
        .I3(\processor/mem_rd_address [4]),
        .I4(\processor/execute/rs2_addr [4]),
        .O(registers_reg_r1_0_31_0_5_i_12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    registers_reg_r1_0_31_0_5_i_13
       (.I0(\processor/execute/rs2_addr [4]),
        .I1(\processor/execute/rs2_addr [1]),
        .I2(\processor/execute/rs2_addr [0]),
        .I3(\processor/execute/rs2_addr [3]),
        .I4(\processor/execute/rs2_addr [2]),
        .O(registers_reg_r1_0_31_0_5_i_13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    registers_reg_r1_0_31_0_5_i_14
       (.I0(\processor/execute/rs1_addr[0]_repN ),
        .I1(\processor/mem_rd_address [0]),
        .I2(\processor/mem_rd_address [1]),
        .I3(\processor/execute/rs1_addr [1]),
        .I4(\processor/mem_rd_address [2]),
        .I5(\processor/execute/rs1_addr [2]),
        .O(registers_reg_r1_0_31_0_5_i_14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE2)) 
    registers_reg_r1_0_31_0_5_i_2
       (.I0(\processor/rs2_address_p [4]),
        .I1(\processor/execute/exception_taken0 ),
        .I2(\processor/id_shamt [4]),
        .O(\processor/rs2_address [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE2)) 
    registers_reg_r1_0_31_0_5_i_3
       (.I0(\processor/rs2_address_p [3]),
        .I1(\processor/execute/exception_taken0 ),
        .I2(\processor/id_shamt [3]),
        .O(\processor/rs2_address [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE2)) 
    registers_reg_r1_0_31_0_5_i_4
       (.I0(\processor/rs2_address_p [2]),
        .I1(\processor/execute/exception_taken0 ),
        .I2(\processor/id_shamt [2]),
        .O(\processor/rs2_address [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE2)) 
    registers_reg_r1_0_31_0_5_i_5
       (.I0(\processor/rs2_address_p [1]),
        .I1(\processor/execute/exception_taken0 ),
        .I2(\processor/id_shamt [1]),
        .O(\processor/rs2_address [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE2)) 
    registers_reg_r1_0_31_0_5_i_6
       (.I0(\processor/rs2_address_p [0]),
        .I1(\processor/execute/exception_taken0 ),
        .I2(\processor/id_shamt [0]),
        .O(\processor/rs2_address [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBBBF0000)) 
    registers_reg_r1_0_31_0_5_i_7
       (.I0(\processor/mem_mem_op [2]),
        .I1(\processor/mem_mem_op [1]),
        .I2(registers_reg_r1_0_31_0_5_i_8_n_0),
        .I3(registers_reg_r1_0_31_0_5_i_9_n_0),
        .I4(\processor/memory/p_1_in ),
        .O(\processor/execute/exception_taken0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000002)) 
    registers_reg_r1_0_31_0_5_i_8
       (.I0(registers_reg_r1_0_31_0_5_i_10_n_0),
        .I1(\processor/execute/alu_x_src [1]),
        .I2(\processor/execute/alu_x_src [0]),
        .I3(\processor/execute/alu_x_src [2]),
        .I4(registers_reg_r1_0_31_0_5_i_11_n_0),
        .O(registers_reg_r1_0_31_0_5_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000002)) 
    registers_reg_r1_0_31_0_5_i_9
       (.I0(registers_reg_r1_0_31_0_5_i_12_n_0),
        .I1(\processor/execute/alu_y_src [2]),
        .I2(\processor/execute/alu_y_src [0]),
        .I3(\processor/execute/alu_y_src [1]),
        .I4(registers_reg_r1_0_31_0_5_i_13_n_0),
        .O(registers_reg_r1_0_31_0_5_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE2)) 
    registers_reg_r2_0_31_0_5_i_1
       (.I0(\processor/rs1_address_p [4]),
        .I1(\processor/execute/exception_taken0 ),
        .I2(\processor/id_rs1_address [4]),
        .O(\processor/rs1_address [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE2)) 
    registers_reg_r2_0_31_0_5_i_2
       (.I0(\processor/rs1_address_p [3]),
        .I1(\processor/execute/exception_taken0 ),
        .I2(\processor/id_rs1_address [3]),
        .O(\processor/rs1_address [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE2)) 
    registers_reg_r2_0_31_0_5_i_3
       (.I0(\processor/rs1_address_p [2]),
        .I1(\processor/execute/exception_taken0 ),
        .I2(\processor/id_rs1_address [2]),
        .O(\processor/rs1_address [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE2)) 
    registers_reg_r2_0_31_0_5_i_4
       (.I0(\processor/rs1_address_p [1]),
        .I1(\processor/execute/exception_taken0 ),
        .I2(\processor/id_rs1_address [1]),
        .O(\processor/rs1_address [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE2)) 
    registers_reg_r2_0_31_0_5_i_5
       (.I0(\processor/rs1_address_p [0]),
        .I1(\processor/execute/exception_taken0 ),
        .I2(\processor/id_rs1_address [0]),
        .O(\processor/rs1_address [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair189" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[0]_i_1 
       (.I0(\processor/wb_rd_data [0]),
        .I1(rs1_data),
        .I2(p_1_out0_in[0]),
        .O(p_1_out2_out[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair180" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[10]_i_1 
       (.I0(\processor/wb_rd_data [10]),
        .I1(rs1_data),
        .I2(p_1_out0_in[10]),
        .O(p_1_out2_out[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair179" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[11]_i_1 
       (.I0(\processor/wb_rd_data [11]),
        .I1(rs1_data),
        .I2(p_1_out0_in[11]),
        .O(p_1_out2_out[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair178" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[12]_i_1 
       (.I0(\processor/wb_rd_data [12]),
        .I1(rs1_data),
        .I2(p_1_out0_in[12]),
        .O(p_1_out2_out[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair177" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[13]_i_1 
       (.I0(\processor/wb_rd_data [13]),
        .I1(rs1_data),
        .I2(p_1_out0_in[13]),
        .O(p_1_out2_out[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair176" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[14]_i_1 
       (.I0(\processor/wb_rd_data [14]),
        .I1(rs1_data),
        .I2(p_1_out0_in[14]),
        .O(p_1_out2_out[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair175" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[15]_i_1 
       (.I0(\processor/wb_rd_data [15]),
        .I1(rs1_data),
        .I2(p_1_out0_in[15]),
        .O(p_1_out2_out[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair174" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[16]_i_1 
       (.I0(\processor/wb_rd_data [16]),
        .I1(rs1_data),
        .I2(p_1_out0_in[16]),
        .O(p_1_out2_out[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair173" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[17]_i_1 
       (.I0(\processor/wb_rd_data [17]),
        .I1(rs1_data),
        .I2(p_1_out0_in[17]),
        .O(p_1_out2_out[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair172" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[18]_i_1 
       (.I0(\processor/wb_rd_data [18]),
        .I1(rs1_data),
        .I2(p_1_out0_in[18]),
        .O(p_1_out2_out[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair171" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[19]_i_1 
       (.I0(\processor/wb_rd_data [19]),
        .I1(rs1_data),
        .I2(p_1_out0_in[19]),
        .O(p_1_out2_out[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair104" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[1]_i_1 
       (.I0(\processor/wb_rd_data [1]),
        .I1(rs1_data),
        .I2(p_1_out0_in[1]),
        .O(p_1_out2_out[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair169" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[20]_i_1 
       (.I0(\processor/wb_rd_data [20]),
        .I1(rs1_data),
        .I2(p_1_out0_in[20]),
        .O(p_1_out2_out[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair168" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[21]_i_1 
       (.I0(\processor/wb_rd_data [21]),
        .I1(rs1_data),
        .I2(p_1_out0_in[21]),
        .O(p_1_out2_out[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair167" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[22]_i_1 
       (.I0(\processor/wb_rd_data [22]),
        .I1(rs1_data),
        .I2(p_1_out0_in[22]),
        .O(p_1_out2_out[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair166" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[23]_i_1 
       (.I0(\processor/wb_rd_data [23]),
        .I1(rs1_data),
        .I2(p_1_out0_in[23]),
        .O(p_1_out2_out[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair165" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[24]_i_1 
       (.I0(\processor/wb_rd_data [24]),
        .I1(rs1_data),
        .I2(p_1_out0_in[24]),
        .O(p_1_out2_out[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair164" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[25]_i_1 
       (.I0(\processor/wb_rd_data [25]),
        .I1(rs1_data),
        .I2(p_1_out0_in[25]),
        .O(p_1_out2_out[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair163" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[26]_i_1 
       (.I0(\processor/wb_rd_data [26]),
        .I1(rs1_data),
        .I2(p_1_out0_in[26]),
        .O(p_1_out2_out[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair162" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[27]_i_1 
       (.I0(\processor/wb_rd_data [27]),
        .I1(rs1_data),
        .I2(p_1_out0_in[27]),
        .O(p_1_out2_out[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair161" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[28]_i_1 
       (.I0(\processor/wb_rd_data [28]),
        .I1(rs1_data),
        .I2(p_1_out0_in[28]),
        .O(p_1_out2_out[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair160" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[29]_i_1 
       (.I0(\processor/wb_rd_data [29]),
        .I1(rs1_data),
        .I2(p_1_out0_in[29]),
        .O(p_1_out2_out[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair188" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[2]_i_1 
       (.I0(\processor/wb_rd_data [2]),
        .I1(rs1_data),
        .I2(p_1_out0_in[2]),
        .O(p_1_out2_out[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair159" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[30]_i_1 
       (.I0(\processor/wb_rd_data [30]),
        .I1(rs1_data),
        .I2(p_1_out0_in[30]),
        .O(p_1_out2_out[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair158" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[31]_i_1 
       (.I0(\processor/wb_rd_data [31]),
        .I1(rs1_data),
        .I2(p_1_out0_in[31]),
        .O(p_1_out2_out[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8200000000008200)) 
    \rs1_data[31]_i_2 
       (.I0(\processor/regfile/p_0_in ),
        .I1(\processor/rs1_address [4]),
        .I2(\processor/wb_rd_address [4]),
        .I3(\rs1_data[31]_i_3_n_0 ),
        .I4(\processor/wb_rd_address [3]),
        .I5(\processor/rs1_address [3]),
        .O(rs1_data));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \rs1_data[31]_i_3 
       (.I0(\processor/rs1_address [0]),
        .I1(\processor/wb_rd_address [0]),
        .I2(\processor/wb_rd_address [2]),
        .I3(\processor/rs1_address [2]),
        .I4(\processor/wb_rd_address [1]),
        .I5(\processor/rs1_address [1]),
        .O(\rs1_data[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair187" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[3]_i_1 
       (.I0(\processor/wb_rd_data [3]),
        .I1(rs1_data),
        .I2(p_1_out0_in[3]),
        .O(p_1_out2_out[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair186" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[4]_i_1 
       (.I0(\processor/wb_rd_data [4]),
        .I1(rs1_data),
        .I2(p_1_out0_in[4]),
        .O(p_1_out2_out[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair185" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[5]_i_1 
       (.I0(\processor/wb_rd_data [5]),
        .I1(rs1_data),
        .I2(p_1_out0_in[5]),
        .O(p_1_out2_out[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair184" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[6]_i_1 
       (.I0(\processor/wb_rd_data [6]),
        .I1(rs1_data),
        .I2(p_1_out0_in[6]),
        .O(p_1_out2_out[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair183" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[7]_i_1 
       (.I0(\processor/wb_rd_data [7]),
        .I1(rs1_data),
        .I2(p_1_out0_in[7]),
        .O(p_1_out2_out[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair182" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[8]_i_1 
       (.I0(\processor/wb_rd_data [8]),
        .I1(rs1_data),
        .I2(p_1_out0_in[8]),
        .O(p_1_out2_out[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair181" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs1_data[9]_i_1 
       (.I0(\processor/wb_rd_data [9]),
        .I1(rs1_data),
        .I2(p_1_out0_in[9]),
        .O(p_1_out2_out[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair189" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[0]_i_1 
       (.I0(\processor/wb_rd_data [0]),
        .I1(rs2_data),
        .I2(p_2_out[0]),
        .O(p_0_out1_out[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair180" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[10]_i_1 
       (.I0(\processor/wb_rd_data [10]),
        .I1(rs2_data),
        .I2(p_2_out[10]),
        .O(p_0_out1_out[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair179" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[11]_i_1 
       (.I0(\processor/wb_rd_data [11]),
        .I1(rs2_data),
        .I2(p_2_out[11]),
        .O(p_0_out1_out[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair178" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[12]_i_1 
       (.I0(\processor/wb_rd_data [12]),
        .I1(rs2_data),
        .I2(p_2_out[12]),
        .O(p_0_out1_out[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair177" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[13]_i_1 
       (.I0(\processor/wb_rd_data [13]),
        .I1(rs2_data),
        .I2(p_2_out[13]),
        .O(p_0_out1_out[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair176" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[14]_i_1 
       (.I0(\processor/wb_rd_data [14]),
        .I1(rs2_data),
        .I2(p_2_out[14]),
        .O(p_0_out1_out[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair175" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[15]_i_1 
       (.I0(\processor/wb_rd_data [15]),
        .I1(rs2_data),
        .I2(p_2_out[15]),
        .O(p_0_out1_out[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair174" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[16]_i_1 
       (.I0(\processor/wb_rd_data [16]),
        .I1(rs2_data),
        .I2(p_2_out[16]),
        .O(p_0_out1_out[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair173" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[17]_i_1 
       (.I0(\processor/wb_rd_data [17]),
        .I1(rs2_data),
        .I2(p_2_out[17]),
        .O(p_0_out1_out[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair172" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[18]_i_1 
       (.I0(\processor/wb_rd_data [18]),
        .I1(rs2_data),
        .I2(p_2_out[18]),
        .O(p_0_out1_out[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair171" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[19]_i_1 
       (.I0(\processor/wb_rd_data [19]),
        .I1(rs2_data),
        .I2(p_2_out[19]),
        .O(p_0_out1_out[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair104" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[1]_i_1 
       (.I0(\processor/wb_rd_data [1]),
        .I1(rs2_data),
        .I2(p_2_out[1]),
        .O(p_0_out1_out[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair169" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[20]_i_1 
       (.I0(\processor/wb_rd_data [20]),
        .I1(rs2_data),
        .I2(p_2_out[20]),
        .O(p_0_out1_out[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair168" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[21]_i_1 
       (.I0(\processor/wb_rd_data [21]),
        .I1(rs2_data),
        .I2(p_2_out[21]),
        .O(p_0_out1_out[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair167" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[22]_i_1 
       (.I0(\processor/wb_rd_data [22]),
        .I1(rs2_data),
        .I2(p_2_out[22]),
        .O(p_0_out1_out[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair166" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[23]_i_1 
       (.I0(\processor/wb_rd_data [23]),
        .I1(rs2_data),
        .I2(p_2_out[23]),
        .O(p_0_out1_out[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair165" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[24]_i_1 
       (.I0(\processor/wb_rd_data [24]),
        .I1(rs2_data),
        .I2(p_2_out[24]),
        .O(p_0_out1_out[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair164" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[25]_i_1 
       (.I0(\processor/wb_rd_data [25]),
        .I1(rs2_data),
        .I2(p_2_out[25]),
        .O(p_0_out1_out[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair163" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[26]_i_1 
       (.I0(\processor/wb_rd_data [26]),
        .I1(rs2_data),
        .I2(p_2_out[26]),
        .O(p_0_out1_out[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair162" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[27]_i_1 
       (.I0(\processor/wb_rd_data [27]),
        .I1(rs2_data),
        .I2(p_2_out[27]),
        .O(p_0_out1_out[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair161" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[28]_i_1 
       (.I0(\processor/wb_rd_data [28]),
        .I1(rs2_data),
        .I2(p_2_out[28]),
        .O(p_0_out1_out[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair160" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[29]_i_1 
       (.I0(\processor/wb_rd_data [29]),
        .I1(rs2_data),
        .I2(p_2_out[29]),
        .O(p_0_out1_out[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair188" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[2]_i_1 
       (.I0(\processor/wb_rd_data [2]),
        .I1(rs2_data),
        .I2(p_2_out[2]),
        .O(p_0_out1_out[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair159" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[30]_i_1 
       (.I0(\processor/wb_rd_data [30]),
        .I1(rs2_data),
        .I2(p_2_out[30]),
        .O(p_0_out1_out[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair158" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[31]_i_1 
       (.I0(\processor/wb_rd_data [31]),
        .I1(rs2_data),
        .I2(p_2_out[31]),
        .O(p_0_out1_out[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8200000000008200)) 
    \rs2_data[31]_i_2 
       (.I0(\processor/regfile/p_0_in ),
        .I1(\processor/rs2_address [4]),
        .I2(\processor/wb_rd_address [4]),
        .I3(\rs2_data[31]_i_3_n_0 ),
        .I4(\processor/wb_rd_address [3]),
        .I5(\processor/rs2_address [3]),
        .O(rs2_data));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \rs2_data[31]_i_3 
       (.I0(\processor/rs2_address [0]),
        .I1(\processor/wb_rd_address [0]),
        .I2(\processor/wb_rd_address [2]),
        .I3(\processor/rs2_address [2]),
        .I4(\processor/wb_rd_address [1]),
        .I5(\processor/rs2_address [1]),
        .O(\rs2_data[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair187" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[3]_i_1 
       (.I0(\processor/wb_rd_data [3]),
        .I1(rs2_data),
        .I2(p_2_out[3]),
        .O(p_0_out1_out[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair186" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[4]_i_1 
       (.I0(\processor/wb_rd_data [4]),
        .I1(rs2_data),
        .I2(p_2_out[4]),
        .O(p_0_out1_out[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair185" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[5]_i_1 
       (.I0(\processor/wb_rd_data [5]),
        .I1(rs2_data),
        .I2(p_2_out[5]),
        .O(p_0_out1_out[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair184" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[6]_i_1 
       (.I0(\processor/wb_rd_data [6]),
        .I1(rs2_data),
        .I2(p_2_out[6]),
        .O(p_0_out1_out[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair183" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[7]_i_1 
       (.I0(\processor/wb_rd_data [7]),
        .I1(rs2_data),
        .I2(p_2_out[7]),
        .O(p_0_out1_out[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair182" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[8]_i_1 
       (.I0(\processor/wb_rd_data [8]),
        .I1(rs2_data),
        .I2(p_2_out[8]),
        .O(p_0_out1_out[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair181" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \rs2_data[9]_i_1 
       (.I0(\processor/wb_rd_data [9]),
        .I1(rs2_data),
        .I2(p_2_out[9]),
        .O(p_0_out1_out[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFABFFFF00A80000)) 
    software_interrupt_i_1
       (.I0(\processor/wb_csr_data [3]),
        .I1(\processor/wb_csr_write [0]),
        .I2(\processor/wb_csr_write [1]),
        .I3(\mtime_compare[31]_i_3_n_0 ),
        .I4(\processor/csr_unit/software_interrupt__5 ),
        .I5(\processor/software_interrupt ),
        .O(software_interrupt_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    software_interrupt_i_2
       (.I0(\processor/wb_csr_address [5]),
        .I1(\processor/wb_csr_address [1]),
        .I2(\processor/wb_csr_address [2]),
        .I3(\processor/wb_csr_address [6]),
        .I4(\processor/wb_csr_address [0]),
        .I5(\mtime_compare[31]_i_4_n_0 ),
        .O(\processor/csr_unit/software_interrupt__5 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair38" *) 
  LUT4 #(
    .INIT(16'h44EC)) 
    \state[0]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[2] ),
        .I2(\icache/state_reg_n_0_[1] ),
        .I3(icache_inputs),
        .O(state));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0200FFFF02000000)) 
    \state[1]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\state[1]_i_2__0_n_0 ),
        .I2(\icache/cl_current_word_reg_n_0_[2] ),
        .I3(\icache/state_reg_n_0_[2] ),
        .I4(\state[1]_i_3__0_n_0 ),
        .I5(\icache/state_reg_n_0_[1] ),
        .O(\state[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2222222222222E22)) 
    \state[1]_i_2 
       (.I0(\processor/dmem_write_req_p ),
        .I1(\processor/memory/p_1_in ),
        .I2(\processor/ex_mem_op [0]),
        .I3(\processor/ex_mem_op [2]),
        .I4(\processor/ex_mem_op [1]),
        .I5(\mem_op[2]_i_5_n_0 ),
        .O(dmem_write_req));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \state[1]_i_2__0 
       (.I0(\icache/cl_current_word_reg_n_0_[1] ),
        .I1(\icache/cl_current_word_reg_n_0_ ),
        .O(\state[1]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000755530002000)) 
    \state[1]_i_3 
       (.I0(\dmem_if/state_reg_n_0_[1] ),
        .I1(\arbiter/state [0]),
        .I2(wb_ack_in),
        .I3(\arbiter/state [1]),
        .I4(\dmem_if/state_reg_n_0_ ),
        .I5(\wb_outputs[adr][31]_i_3_n_0 ),
        .O(\state[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFD303D)) 
    \state[1]_i_3__0 
       (.I0(\icache/cache_hit ),
        .I1(\icache/state_reg_n_0_ ),
        .I2(\icache/state_reg_n_0_[2] ),
        .I3(\icache/state_reg_n_0_[1] ),
        .I4(icache_inputs),
        .O(\state[1]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00F1C0F1)) 
    \state[2]_i_1 
       (.I0(\icache/cache_hit ),
        .I1(\icache/state_reg_n_0_ ),
        .I2(\icache/state_reg_n_0_[2] ),
        .I3(\icache/state_reg_n_0_[1] ),
        .I4(icache_inputs),
        .O(\state[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5555FFFF00008000)) 
    store_cache_line_i_1
       (.I0(\icache/state_reg_n_0_[2] ),
        .I1(\icache/state_reg_n_0_ ),
        .I2(\icache/store_cache_line__1 ),
        .I3(icache_inputs),
        .I4(\icache/state_reg_n_0_[1] ),
        .I5(\icache/store_cache_line_reg_n_0 ),
        .O(store_cache_line_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    store_cache_line_i_2
       (.I0(\icache/cl_current_word_reg_n_0_[2] ),
        .I1(\icache/cl_current_word_reg_n_0_ ),
        .I2(\icache/cl_current_word_reg_n_0_[1] ),
        .O(\icache/store_cache_line__1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    tag_memory_reg_0_63_0_2_i_1
       (.I0(reset),
        .I1(\icache/store_cache_line_reg_n_0 ),
        .I2(\icache/cl_load_address [10]),
        .O(tag_memory_reg_0_63_0_2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    tag_memory_reg_0_63_0_2_i_10
       (.I0(\processor/mem_csr_data [4]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [4]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [4]),
        .O(\processor/exception_target [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    tag_memory_reg_0_63_0_2_i_11
       (.I0(\pc[4]_i_2_n_0 ),
        .I1(\mem_op[2]_i_4_n_0 ),
        .I2(\pc_reg[4]_i_3_n_4 ),
        .O(tag_memory_reg_0_63_0_2_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    tag_memory_reg_0_63_0_2_i_12
       (.I0(\processor/mem_csr_data [7]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [7]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [7]),
        .O(\processor/execute/mtvec_forwarded [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    tag_memory_reg_0_63_0_2_i_13
       (.I0(\processor/mem_csr_data [6]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [6]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [6]),
        .O(\processor/execute/mtvec_forwarded [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    tag_memory_reg_0_63_0_2_i_14
       (.I0(\processor/mem_csr_data [8]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [8]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [8]),
        .O(\processor/execute/mtvec_forwarded [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h001DFF1D)) 
    tag_memory_reg_0_63_0_2_i_15
       (.I0(\processor/execute/mtvec [7]),
        .I1(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I2(\processor/wb_csr_data [7]),
        .I3(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I4(\processor/mem_csr_data [7]),
        .O(tag_memory_reg_0_63_0_2_i_15_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h001DFF1D)) 
    tag_memory_reg_0_63_0_2_i_16
       (.I0(\processor/execute/mtvec [6]),
        .I1(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I2(\processor/wb_csr_data [6]),
        .I3(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I4(\processor/mem_csr_data [6]),
        .O(tag_memory_reg_0_63_0_2_i_16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    tag_memory_reg_0_63_0_2_i_17
       (.I0(\processor/mem_csr_data [5]),
        .I1(tag_memory_reg_0_63_0_2_i_18_n_0),
        .I2(\processor/wb_csr_data [5]),
        .I3(tag_memory_reg_0_63_0_2_i_19_n_0),
        .I4(\processor/execute/mtvec [5]),
        .O(\processor/execute/mtvec_forwarded [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    tag_memory_reg_0_63_0_2_i_18
       (.I0(tag_memory_reg_0_63_0_2_i_20_n_0),
        .I1(\processor/mem_csr_address [7]),
        .I2(\processor/mem_csr_address [1]),
        .I3(\processor/mem_csr_address [10]),
        .I4(\processor/mem_csr_address [2]),
        .I5(\processor/mem_csr_address [0]),
        .O(tag_memory_reg_0_63_0_2_i_18_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000200000000000)) 
    tag_memory_reg_0_63_0_2_i_19
       (.I0(tag_memory_reg_0_63_0_2_i_21_n_0),
        .I1(\processor/wb_csr_address [10]),
        .I2(\processor/wb_csr_address [9]),
        .I3(\processor/wb_csr_address [8]),
        .I4(\processor/wb_csr_address [4]),
        .I5(\processor/csr_unit/tohost_data1__0 ),
        .O(tag_memory_reg_0_63_0_2_i_19_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    tag_memory_reg_0_63_0_2_i_2
       (.I0(pc[9]),
        .I1(pc_next[9]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0002000200020000)) 
    tag_memory_reg_0_63_0_2_i_20
       (.I0(\exception_context_out[ie1]_i_7_n_0 ),
        .I1(\processor/mem_csr_address [4]),
        .I2(\processor/mem_csr_address [11]),
        .I3(\processor/mem_csr_address [3]),
        .I4(\processor/mem_csr_write [0]),
        .I5(\processor/mem_csr_write [1]),
        .O(tag_memory_reg_0_63_0_2_i_20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    tag_memory_reg_0_63_0_2_i_21
       (.I0(tag_memory_reg_0_63_0_2_i_22_n_0),
        .I1(\processor/wb_csr_address [0]),
        .I2(\processor/wb_csr_address [2]),
        .I3(\processor/wb_csr_address [1]),
        .I4(\processor/wb_csr_address [7]),
        .I5(tag_memory_reg_0_63_0_2_i_23_n_0),
        .O(tag_memory_reg_0_63_0_2_i_21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    tag_memory_reg_0_63_0_2_i_22
       (.I0(\processor/wb_csr_address [5]),
        .I1(\processor/wb_csr_address [6]),
        .O(tag_memory_reg_0_63_0_2_i_22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    tag_memory_reg_0_63_0_2_i_23
       (.I0(\processor/wb_csr_address [3]),
        .I1(\processor/wb_csr_address [11]),
        .O(tag_memory_reg_0_63_0_2_i_23_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    tag_memory_reg_0_63_0_2_i_3
       (.I0(pc[8]),
        .I1(pc_next[8]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    tag_memory_reg_0_63_0_2_i_4
       (.I0(pc[7]),
        .I1(pc_next[7]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    tag_memory_reg_0_63_0_2_i_5
       (.I0(pc[6]),
        .I1(pc_next[6]),
        .I2(\processor/fetch/cancel_fetch ),
        .O(imem_address[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACCF0)) 
    tag_memory_reg_0_63_0_2_i_6
       (.I0(pc[5]),
        .I1(\processor/exception_target [5]),
        .I2(tag_memory_reg_0_63_0_2_i_9_n_0),
        .I3(\mem_op[2]_i_5_n_0 ),
        .I4(\processor/fetch/cancel_fetch ),
        .O(imem_address[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAACCF0)) 
    tag_memory_reg_0_63_0_2_i_7
       (.I0(pc[4]),
        .I1(\processor/exception_target [4]),
        .I2(tag_memory_reg_0_63_0_2_i_11_n_0),
        .I3(\mem_op[2]_i_5_n_0 ),
        .I4(\processor/fetch/cancel_fetch ),
        .O(imem_address[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 tag_memory_reg_0_63_0_2_i_8
       (.CI(\<const0>__0__0 ),
        .CO({tag_memory_reg_0_63_0_2_i_8_n_0,tag_memory_reg_0_63_0_2_i_8_n_1,tag_memory_reg_0_63_0_2_i_8_n_2,tag_memory_reg_0_63_0_2_i_8_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\processor/execute/mtvec_forwarded [7:6],\<const0>__0__0 }),
        .O(\processor/exception_target [8:5]),
        .S({\processor/execute/mtvec_forwarded [8],tag_memory_reg_0_63_0_2_i_15_n_0,tag_memory_reg_0_63_0_2_i_16_n_0,\processor/execute/mtvec_forwarded [5]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    tag_memory_reg_0_63_0_2_i_9
       (.I0(\pc[5]_i_2_n_0 ),
        .I1(\mem_op[2]_i_4_n_0 ),
        .I2(\pc_reg[8]_i_3_n_7 ),
        .O(tag_memory_reg_0_63_0_2_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    tag_memory_reg_64_127_0_2_i_1
       (.I0(reset),
        .I1(\icache/store_cache_line_reg_n_0 ),
        .I2(\icache/cl_load_address [10]),
        .O(tag_memory_reg_64_127_0_2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    timer_interrupt0_inferred__0_carry__0_i_1
       (.I0(\processor/csr_unit/counter_mtime_reg [21]),
        .I1(mtime_compare[21]),
        .I2(mtime_compare[23]),
        .I3(\processor/csr_unit/counter_mtime_reg [23]),
        .I4(mtime_compare[22]),
        .I5(\processor/csr_unit/counter_mtime_reg [22]),
        .O(timer_interrupt0_inferred__0_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    timer_interrupt0_inferred__0_carry__0_i_2
       (.I0(\processor/csr_unit/counter_mtime_reg [18]),
        .I1(mtime_compare[18]),
        .I2(mtime_compare[20]),
        .I3(\processor/csr_unit/counter_mtime_reg [20]),
        .I4(mtime_compare[19]),
        .I5(\processor/csr_unit/counter_mtime_reg [19]),
        .O(timer_interrupt0_inferred__0_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    timer_interrupt0_inferred__0_carry__0_i_3
       (.I0(\processor/csr_unit/counter_mtime_reg [15]),
        .I1(mtime_compare[15]),
        .I2(mtime_compare[17]),
        .I3(\processor/csr_unit/counter_mtime_reg [17]),
        .I4(mtime_compare[16]),
        .I5(\processor/csr_unit/counter_mtime_reg [16]),
        .O(timer_interrupt0_inferred__0_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    timer_interrupt0_inferred__0_carry__0_i_4
       (.I0(\processor/csr_unit/counter_mtime_reg [12]),
        .I1(mtime_compare[12]),
        .I2(mtime_compare[14]),
        .I3(\processor/csr_unit/counter_mtime_reg [14]),
        .I4(mtime_compare[13]),
        .I5(\processor/csr_unit/counter_mtime_reg [13]),
        .O(timer_interrupt0_inferred__0_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    timer_interrupt0_inferred__0_carry__1_i_1
       (.I0(\processor/csr_unit/counter_mtime_reg [30]),
        .I1(mtime_compare[30]),
        .I2(\processor/csr_unit/counter_mtime_reg [31]),
        .I3(mtime_compare[31]),
        .O(timer_interrupt0_inferred__0_carry__1_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    timer_interrupt0_inferred__0_carry__1_i_2
       (.I0(\processor/csr_unit/counter_mtime_reg [27]),
        .I1(mtime_compare[27]),
        .I2(mtime_compare[29]),
        .I3(\processor/csr_unit/counter_mtime_reg [29]),
        .I4(mtime_compare[28]),
        .I5(\processor/csr_unit/counter_mtime_reg [28]),
        .O(timer_interrupt0_inferred__0_carry__1_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    timer_interrupt0_inferred__0_carry__1_i_3
       (.I0(\processor/csr_unit/counter_mtime_reg [24]),
        .I1(mtime_compare[24]),
        .I2(mtime_compare[26]),
        .I3(\processor/csr_unit/counter_mtime_reg [26]),
        .I4(mtime_compare[25]),
        .I5(\processor/csr_unit/counter_mtime_reg [25]),
        .O(timer_interrupt0_inferred__0_carry__1_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    timer_interrupt0_inferred__0_carry_i_1
       (.I0(\processor/csr_unit/counter_mtime_reg [9]),
        .I1(mtime_compare[9]),
        .I2(mtime_compare[11]),
        .I3(\processor/csr_unit/counter_mtime_reg [11]),
        .I4(mtime_compare[10]),
        .I5(\processor/csr_unit/counter_mtime_reg [10]),
        .O(timer_interrupt0_inferred__0_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    timer_interrupt0_inferred__0_carry_i_2
       (.I0(\processor/csr_unit/counter_mtime_reg [6]),
        .I1(mtime_compare[6]),
        .I2(mtime_compare[8]),
        .I3(\processor/csr_unit/counter_mtime_reg [8]),
        .I4(mtime_compare[7]),
        .I5(\processor/csr_unit/counter_mtime_reg [7]),
        .O(timer_interrupt0_inferred__0_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    timer_interrupt0_inferred__0_carry_i_3
       (.I0(\processor/csr_unit/counter_mtime_reg [3]),
        .I1(mtime_compare[3]),
        .I2(mtime_compare[5]),
        .I3(\processor/csr_unit/counter_mtime_reg [5]),
        .I4(mtime_compare[4]),
        .I5(\processor/csr_unit/counter_mtime_reg [4]),
        .O(timer_interrupt0_inferred__0_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    timer_interrupt0_inferred__0_carry_i_4
       (.I0(\processor/csr_unit/counter_mtime_reg [0]),
        .I1(mtime_compare[0]),
        .I2(mtime_compare[2]),
        .I3(\processor/csr_unit/counter_mtime_reg [2]),
        .I4(mtime_compare[1]),
        .I5(\processor/csr_unit/counter_mtime_reg [1]),
        .O(timer_interrupt0_inferred__0_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h000E)) 
    timer_interrupt_i_1
       (.I0(\processor/timer_interrupt ),
        .I1(\processor/csr_unit/timer_interrupt0_inferred__0_carry__1_n_1 ),
        .I2(\processor/csr_unit/timer_interrupt0__8 ),
        .I3(reset),
        .O(timer_interrupt_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    timer_interrupt_i_2
       (.I0(timer_interrupt_i_3_n_0),
        .I1(timer_interrupt_i_4_n_0),
        .I2(\processor/wb_csr_address [6]),
        .I3(\processor/wb_csr_address [7]),
        .I4(\processor/wb_csr_address [4]),
        .I5(\processor/wb_csr_address [2]),
        .O(\processor/csr_unit/timer_interrupt0__8 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF1)) 
    timer_interrupt_i_3
       (.I0(\processor/wb_csr_write [0]),
        .I1(\processor/wb_csr_write [1]),
        .I2(\processor/wb_csr_address [3]),
        .I3(\processor/wb_csr_address [1]),
        .I4(\processor/wb_csr_address [11]),
        .I5(\processor/wb_csr_address [10]),
        .O(timer_interrupt_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    timer_interrupt_i_4
       (.I0(\processor/wb_csr_address [5]),
        .I1(\processor/wb_csr_address [9]),
        .I2(\processor/wb_csr_address [0]),
        .I3(\processor/wb_csr_address [8]),
        .O(timer_interrupt_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \tohost_data[31]_i_1 
       (.I0(\processor/wb_csr_address [11]),
        .I1(\processor/wb_csr_address [3]),
        .I2(\processor/wb_csr_address [1]),
        .I3(\processor/wb_csr_address [0]),
        .I4(\processor/csr_unit/tohost_data1__0 ),
        .I5(\tohost_data[31]_i_3_n_0 ),
        .O(\processor/csr_unit/tohost_data0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \tohost_data[31]_i_2 
       (.I0(\processor/wb_csr_write [1]),
        .I1(\processor/wb_csr_write [0]),
        .O(\processor/csr_unit/tohost_data1__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFEFFFFFFFFFFFF)) 
    \tohost_data[31]_i_3 
       (.I0(\processor/wb_csr_address [5]),
        .I1(\processor/wb_csr_address [4]),
        .I2(\tohost_data[31]_i_4_n_0 ),
        .I3(\tohost_data[31]_i_5_n_0 ),
        .I4(\processor/wb_csr_address [10]),
        .I5(\processor/wb_csr_address [7]),
        .O(\tohost_data[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \tohost_data[31]_i_4 
       (.I0(\processor/wb_csr_address [2]),
        .I1(\processor/wb_csr_address [6]),
        .O(\tohost_data[31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \tohost_data[31]_i_5 
       (.I0(\processor/wb_csr_address [8]),
        .I1(\processor/wb_csr_address [9]),
        .O(\tohost_data[31]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[0]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[112]_i_2_n_0 ),
        .I3(\valid[15]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [0]),
        .O(valid));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[100]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[116]_i_2_n_0 ),
        .I3(\valid[111]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [100]),
        .O(\valid[100]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[101]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[117]_i_2_n_0 ),
        .I3(\valid[111]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [101]),
        .O(\valid[101]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[102]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[118]_i_2_n_0 ),
        .I3(\valid[111]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [102]),
        .O(\valid[102]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[103]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[119]_i_2_n_0 ),
        .I3(\valid[111]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [103]),
        .O(\valid[103]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[104]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[120]_i_2_n_0 ),
        .I3(\valid[111]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [104]),
        .O(\valid[104]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[105]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[121]_i_2_n_0 ),
        .I3(\valid[111]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [105]),
        .O(\valid[105]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[106]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[122]_i_2_n_0 ),
        .I3(\valid[111]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [106]),
        .O(\valid[106]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[107]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[123]_i_2_n_0 ),
        .I3(\valid[111]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [107]),
        .O(\valid[107]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[108]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[124]_i_2_n_0 ),
        .I3(\valid[111]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [108]),
        .O(\valid[108]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[109]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[125]_i_2_n_0 ),
        .I3(\valid[111]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [109]),
        .O(\valid[109]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[10]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[122]_i_2_n_0 ),
        .I3(\valid[15]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [10]),
        .O(\valid[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[110]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[126]_i_2_n_0 ),
        .I3(\valid[111]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [110]),
        .O(\valid[110]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[111]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[127]_i_2_n_0 ),
        .I3(\valid[111]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [111]),
        .O(\valid[111]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hDF)) 
    \valid[111]_i_2 
       (.I0(\icache/cl_load_address [10]),
        .I1(\icache/cl_load_address [8]),
        .I2(\icache/cl_load_address [9]),
        .O(\valid[111]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[112]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[112]_i_2_n_0 ),
        .I3(\valid[127]_i_3_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [112]),
        .O(\valid[112]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \valid[112]_i_2 
       (.I0(\icache/cl_load_address [6]),
        .I1(\icache/cl_load_address [7]),
        .I2(\icache/cl_load_address [4]),
        .I3(\icache/cl_load_address [5]),
        .O(\valid[112]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[113]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[113]_i_2_n_0 ),
        .I3(\valid[127]_i_3_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [113]),
        .O(\valid[113]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFEFF)) 
    \valid[113]_i_2 
       (.I0(\icache/cl_load_address [6]),
        .I1(\icache/cl_load_address [7]),
        .I2(\icache/cl_load_address [5]),
        .I3(\icache/cl_load_address [4]),
        .O(\valid[113]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[114]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[114]_i_2_n_0 ),
        .I3(\valid[127]_i_3_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [114]),
        .O(\valid[114]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFEFF)) 
    \valid[114]_i_2 
       (.I0(\icache/cl_load_address [6]),
        .I1(\icache/cl_load_address [7]),
        .I2(\icache/cl_load_address [4]),
        .I3(\icache/cl_load_address [5]),
        .O(\valid[114]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[115]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[115]_i_2_n_0 ),
        .I3(\valid[127]_i_3_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [115]),
        .O(\valid[115]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEFFF)) 
    \valid[115]_i_2 
       (.I0(\icache/cl_load_address [6]),
        .I1(\icache/cl_load_address [7]),
        .I2(\icache/cl_load_address [4]),
        .I3(\icache/cl_load_address [5]),
        .O(\valid[115]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[116]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[116]_i_2_n_0 ),
        .I3(\valid[127]_i_3_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [116]),
        .O(\valid[116]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFB)) 
    \valid[116]_i_2 
       (.I0(\icache/cl_load_address [7]),
        .I1(\icache/cl_load_address [6]),
        .I2(\icache/cl_load_address [4]),
        .I3(\icache/cl_load_address [5]),
        .O(\valid[116]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[117]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[117]_i_2_n_0 ),
        .I3(\valid[127]_i_3_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [117]),
        .O(\valid[117]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFBFF)) 
    \valid[117]_i_2 
       (.I0(\icache/cl_load_address [7]),
        .I1(\icache/cl_load_address [6]),
        .I2(\icache/cl_load_address [5]),
        .I3(\icache/cl_load_address [4]),
        .O(\valid[117]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[118]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[118]_i_2_n_0 ),
        .I3(\valid[127]_i_3_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [118]),
        .O(\valid[118]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFBFF)) 
    \valid[118]_i_2 
       (.I0(\icache/cl_load_address [7]),
        .I1(\icache/cl_load_address [6]),
        .I2(\icache/cl_load_address [4]),
        .I3(\icache/cl_load_address [5]),
        .O(\valid[118]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[119]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[119]_i_2_n_0 ),
        .I3(\valid[127]_i_3_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [119]),
        .O(\valid[119]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBFFF)) 
    \valid[119]_i_2 
       (.I0(\icache/cl_load_address [7]),
        .I1(\icache/cl_load_address [6]),
        .I2(\icache/cl_load_address [4]),
        .I3(\icache/cl_load_address [5]),
        .O(\valid[119]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[11]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[123]_i_2_n_0 ),
        .I3(\valid[15]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [11]),
        .O(\valid[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[120]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[120]_i_2_n_0 ),
        .I3(\valid[127]_i_3_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [120]),
        .O(\valid[120]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFB)) 
    \valid[120]_i_2 
       (.I0(\icache/cl_load_address [6]),
        .I1(\icache/cl_load_address [7]),
        .I2(\icache/cl_load_address [4]),
        .I3(\icache/cl_load_address [5]),
        .O(\valid[120]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[121]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[121]_i_2_n_0 ),
        .I3(\valid[127]_i_3_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [121]),
        .O(\valid[121]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFBFF)) 
    \valid[121]_i_2 
       (.I0(\icache/cl_load_address [6]),
        .I1(\icache/cl_load_address [7]),
        .I2(\icache/cl_load_address [5]),
        .I3(\icache/cl_load_address [4]),
        .O(\valid[121]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[122]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[122]_i_2_n_0 ),
        .I3(\valid[127]_i_3_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [122]),
        .O(\valid[122]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFBFF)) 
    \valid[122]_i_2 
       (.I0(\icache/cl_load_address [6]),
        .I1(\icache/cl_load_address [7]),
        .I2(\icache/cl_load_address [4]),
        .I3(\icache/cl_load_address [5]),
        .O(\valid[122]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[123]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[123]_i_2_n_0 ),
        .I3(\valid[127]_i_3_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [123]),
        .O(\valid[123]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBFFF)) 
    \valid[123]_i_2 
       (.I0(\icache/cl_load_address [6]),
        .I1(\icache/cl_load_address [7]),
        .I2(\icache/cl_load_address [4]),
        .I3(\icache/cl_load_address [5]),
        .O(\valid[123]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[124]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[124]_i_2_n_0 ),
        .I3(\valid[127]_i_3_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [124]),
        .O(\valid[124]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFF7)) 
    \valid[124]_i_2 
       (.I0(\icache/cl_load_address [6]),
        .I1(\icache/cl_load_address [7]),
        .I2(\icache/cl_load_address [4]),
        .I3(\icache/cl_load_address [5]),
        .O(\valid[124]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[125]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[125]_i_2_n_0 ),
        .I3(\valid[127]_i_3_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [125]),
        .O(\valid[125]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF7FF)) 
    \valid[125]_i_2 
       (.I0(\icache/cl_load_address [6]),
        .I1(\icache/cl_load_address [7]),
        .I2(\icache/cl_load_address [5]),
        .I3(\icache/cl_load_address [4]),
        .O(\valid[125]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[126]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[126]_i_2_n_0 ),
        .I3(\valid[127]_i_3_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [126]),
        .O(\valid[126]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF7FF)) 
    \valid[126]_i_2 
       (.I0(\icache/cl_load_address [6]),
        .I1(\icache/cl_load_address [7]),
        .I2(\icache/cl_load_address [4]),
        .I3(\icache/cl_load_address [5]),
        .O(\valid[126]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[127]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[127]_i_2_n_0 ),
        .I3(\valid[127]_i_3_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [127]),
        .O(\valid[127]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    \valid[127]_i_2 
       (.I0(\icache/cl_load_address [6]),
        .I1(\icache/cl_load_address [7]),
        .I2(\icache/cl_load_address [4]),
        .I3(\icache/cl_load_address [5]),
        .O(\valid[127]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h7F)) 
    \valid[127]_i_3 
       (.I0(\icache/cl_load_address [10]),
        .I1(\icache/cl_load_address [8]),
        .I2(\icache/cl_load_address [9]),
        .O(\valid[127]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[12]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[124]_i_2_n_0 ),
        .I3(\valid[15]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [12]),
        .O(\valid[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[13]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[125]_i_2_n_0 ),
        .I3(\valid[15]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [13]),
        .O(\valid[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[14]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[126]_i_2_n_0 ),
        .I3(\valid[15]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [14]),
        .O(\valid[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[15]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[127]_i_2_n_0 ),
        .I3(\valid[15]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [15]),
        .O(\valid[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \valid[15]_i_2 
       (.I0(\icache/cl_load_address [10]),
        .I1(\icache/cl_load_address [8]),
        .I2(\icache/cl_load_address [9]),
        .O(\valid[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[16]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[112]_i_2_n_0 ),
        .I3(\valid[31]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [16]),
        .O(\valid[16]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[17]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[113]_i_2_n_0 ),
        .I3(\valid[31]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [17]),
        .O(\valid[17]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[18]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[114]_i_2_n_0 ),
        .I3(\valid[31]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [18]),
        .O(\valid[18]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[19]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[115]_i_2_n_0 ),
        .I3(\valid[31]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [19]),
        .O(\valid[19]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[1]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[113]_i_2_n_0 ),
        .I3(\valid[15]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [1]),
        .O(\valid[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[20]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[116]_i_2_n_0 ),
        .I3(\valid[31]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [20]),
        .O(\valid[20]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[21]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[117]_i_2_n_0 ),
        .I3(\valid[31]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [21]),
        .O(\valid[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[22]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[118]_i_2_n_0 ),
        .I3(\valid[31]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [22]),
        .O(\valid[22]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[23]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[119]_i_2_n_0 ),
        .I3(\valid[31]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [23]),
        .O(\valid[23]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[24]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[120]_i_2_n_0 ),
        .I3(\valid[31]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [24]),
        .O(\valid[24]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[25]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[121]_i_2_n_0 ),
        .I3(\valid[31]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [25]),
        .O(\valid[25]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[26]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[122]_i_2_n_0 ),
        .I3(\valid[31]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [26]),
        .O(\valid[26]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[27]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[123]_i_2_n_0 ),
        .I3(\valid[31]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [27]),
        .O(\valid[27]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[28]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[124]_i_2_n_0 ),
        .I3(\valid[31]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [28]),
        .O(\valid[28]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[29]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[125]_i_2_n_0 ),
        .I3(\valid[31]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [29]),
        .O(\valid[29]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[2]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[114]_i_2_n_0 ),
        .I3(\valid[15]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [2]),
        .O(\valid[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[30]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[126]_i_2_n_0 ),
        .I3(\valid[31]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [30]),
        .O(\valid[30]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[31]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[127]_i_2_n_0 ),
        .I3(\valid[31]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [31]),
        .O(\valid[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEF)) 
    \valid[31]_i_2 
       (.I0(\icache/cl_load_address [10]),
        .I1(\icache/cl_load_address [9]),
        .I2(\icache/cl_load_address [8]),
        .O(\valid[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[32]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[112]_i_2_n_0 ),
        .I3(\valid[47]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [32]),
        .O(\valid[32]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[33]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[113]_i_2_n_0 ),
        .I3(\valid[47]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [33]),
        .O(\valid[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[34]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[114]_i_2_n_0 ),
        .I3(\valid[47]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [34]),
        .O(\valid[34]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[35]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[115]_i_2_n_0 ),
        .I3(\valid[47]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [35]),
        .O(\valid[35]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[36]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[116]_i_2_n_0 ),
        .I3(\valid[47]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [36]),
        .O(\valid[36]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[37]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[117]_i_2_n_0 ),
        .I3(\valid[47]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [37]),
        .O(\valid[37]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[38]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[118]_i_2_n_0 ),
        .I3(\valid[47]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [38]),
        .O(\valid[38]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[39]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[119]_i_2_n_0 ),
        .I3(\valid[47]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [39]),
        .O(\valid[39]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[3]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[115]_i_2_n_0 ),
        .I3(\valid[15]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [3]),
        .O(\valid[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[40]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[120]_i_2_n_0 ),
        .I3(\valid[47]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [40]),
        .O(\valid[40]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[41]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[121]_i_2_n_0 ),
        .I3(\valid[47]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [41]),
        .O(\valid[41]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[42]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[122]_i_2_n_0 ),
        .I3(\valid[47]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [42]),
        .O(\valid[42]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[43]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[123]_i_2_n_0 ),
        .I3(\valid[47]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [43]),
        .O(\valid[43]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[44]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[124]_i_2_n_0 ),
        .I3(\valid[47]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [44]),
        .O(\valid[44]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[45]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[125]_i_2_n_0 ),
        .I3(\valid[47]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [45]),
        .O(\valid[45]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[46]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[126]_i_2_n_0 ),
        .I3(\valid[47]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [46]),
        .O(\valid[46]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[47]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[127]_i_2_n_0 ),
        .I3(\valid[47]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [47]),
        .O(\valid[47]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEF)) 
    \valid[47]_i_2 
       (.I0(\icache/cl_load_address [10]),
        .I1(\icache/cl_load_address [8]),
        .I2(\icache/cl_load_address [9]),
        .O(\valid[47]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[48]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[112]_i_2_n_0 ),
        .I3(\valid[63]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [48]),
        .O(\valid[48]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[49]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[113]_i_2_n_0 ),
        .I3(\valid[63]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [49]),
        .O(\valid[49]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[4]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[116]_i_2_n_0 ),
        .I3(\valid[15]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [4]),
        .O(\valid[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[50]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[114]_i_2_n_0 ),
        .I3(\valid[63]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [50]),
        .O(\valid[50]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[51]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[115]_i_2_n_0 ),
        .I3(\valid[63]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [51]),
        .O(\valid[51]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[52]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[116]_i_2_n_0 ),
        .I3(\valid[63]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [52]),
        .O(\valid[52]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[53]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[117]_i_2_n_0 ),
        .I3(\valid[63]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [53]),
        .O(\valid[53]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[54]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[118]_i_2_n_0 ),
        .I3(\valid[63]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [54]),
        .O(\valid[54]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[55]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[119]_i_2_n_0 ),
        .I3(\valid[63]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [55]),
        .O(\valid[55]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[56]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[120]_i_2_n_0 ),
        .I3(\valid[63]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [56]),
        .O(\valid[56]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[57]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[121]_i_2_n_0 ),
        .I3(\valid[63]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [57]),
        .O(\valid[57]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[58]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[122]_i_2_n_0 ),
        .I3(\valid[63]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [58]),
        .O(\valid[58]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[59]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[123]_i_2_n_0 ),
        .I3(\valid[63]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [59]),
        .O(\valid[59]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[5]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[117]_i_2_n_0 ),
        .I3(\valid[15]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [5]),
        .O(\valid[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[60]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[124]_i_2_n_0 ),
        .I3(\valid[63]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [60]),
        .O(\valid[60]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[61]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[125]_i_2_n_0 ),
        .I3(\valid[63]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [61]),
        .O(\valid[61]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[62]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[126]_i_2_n_0 ),
        .I3(\valid[63]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [62]),
        .O(\valid[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[63]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[127]_i_2_n_0 ),
        .I3(\valid[63]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [63]),
        .O(\valid[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \valid[63]_i_2 
       (.I0(\icache/cl_load_address [10]),
        .I1(\icache/cl_load_address [8]),
        .I2(\icache/cl_load_address [9]),
        .O(\valid[63]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[64]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[112]_i_2_n_0 ),
        .I3(\valid[79]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [64]),
        .O(\valid[64]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[65]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[113]_i_2_n_0 ),
        .I3(\valid[79]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [65]),
        .O(\valid[65]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[66]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[114]_i_2_n_0 ),
        .I3(\valid[79]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [66]),
        .O(\valid[66]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[67]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[115]_i_2_n_0 ),
        .I3(\valid[79]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [67]),
        .O(\valid[67]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[68]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[116]_i_2_n_0 ),
        .I3(\valid[79]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [68]),
        .O(\valid[68]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[69]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[117]_i_2_n_0 ),
        .I3(\valid[79]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [69]),
        .O(\valid[69]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[6]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[118]_i_2_n_0 ),
        .I3(\valid[15]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [6]),
        .O(\valid[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[70]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[118]_i_2_n_0 ),
        .I3(\valid[79]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [70]),
        .O(\valid[70]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[71]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[119]_i_2_n_0 ),
        .I3(\valid[79]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [71]),
        .O(\valid[71]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[72]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[120]_i_2_n_0 ),
        .I3(\valid[79]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [72]),
        .O(\valid[72]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[73]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[121]_i_2_n_0 ),
        .I3(\valid[79]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [73]),
        .O(\valid[73]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[74]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[122]_i_2_n_0 ),
        .I3(\valid[79]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [74]),
        .O(\valid[74]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[75]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[123]_i_2_n_0 ),
        .I3(\valid[79]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [75]),
        .O(\valid[75]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[76]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[124]_i_2_n_0 ),
        .I3(\valid[79]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [76]),
        .O(\valid[76]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[77]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[125]_i_2_n_0 ),
        .I3(\valid[79]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [77]),
        .O(\valid[77]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[78]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[126]_i_2_n_0 ),
        .I3(\valid[79]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [78]),
        .O(\valid[78]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[79]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[127]_i_2_n_0 ),
        .I3(\valid[79]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [79]),
        .O(\valid[79]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFD)) 
    \valid[79]_i_2 
       (.I0(\icache/cl_load_address [10]),
        .I1(\icache/cl_load_address [8]),
        .I2(\icache/cl_load_address [9]),
        .O(\valid[79]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[7]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[119]_i_2_n_0 ),
        .I3(\valid[15]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [7]),
        .O(\valid[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[80]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[112]_i_2_n_0 ),
        .I3(\valid[95]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [80]),
        .O(\valid[80]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[81]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[113]_i_2_n_0 ),
        .I3(\valid[95]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [81]),
        .O(\valid[81]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[82]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[114]_i_2_n_0 ),
        .I3(\valid[95]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [82]),
        .O(\valid[82]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[83]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[115]_i_2_n_0 ),
        .I3(\valid[95]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [83]),
        .O(\valid[83]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[84]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[116]_i_2_n_0 ),
        .I3(\valid[95]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [84]),
        .O(\valid[84]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[85]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[117]_i_2_n_0 ),
        .I3(\valid[95]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [85]),
        .O(\valid[85]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[86]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[118]_i_2_n_0 ),
        .I3(\valid[95]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [86]),
        .O(\valid[86]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[87]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[119]_i_2_n_0 ),
        .I3(\valid[95]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [87]),
        .O(\valid[87]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[88]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[120]_i_2_n_0 ),
        .I3(\valid[95]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [88]),
        .O(\valid[88]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[89]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[121]_i_2_n_0 ),
        .I3(\valid[95]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [89]),
        .O(\valid[89]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[8]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[120]_i_2_n_0 ),
        .I3(\valid[15]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [8]),
        .O(\valid[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[90]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[122]_i_2_n_0 ),
        .I3(\valid[95]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [90]),
        .O(\valid[90]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[91]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[123]_i_2_n_0 ),
        .I3(\valid[95]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [91]),
        .O(\valid[91]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[92]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[124]_i_2_n_0 ),
        .I3(\valid[95]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [92]),
        .O(\valid[92]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[93]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[125]_i_2_n_0 ),
        .I3(\valid[95]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [93]),
        .O(\valid[93]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[94]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[126]_i_2_n_0 ),
        .I3(\valid[95]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [94]),
        .O(\valid[94]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[95]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[127]_i_2_n_0 ),
        .I3(\valid[95]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [95]),
        .O(\valid[95]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hDF)) 
    \valid[95]_i_2 
       (.I0(\icache/cl_load_address [10]),
        .I1(\icache/cl_load_address [9]),
        .I2(\icache/cl_load_address [8]),
        .O(\valid[95]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[96]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[112]_i_2_n_0 ),
        .I3(\valid[111]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [96]),
        .O(\valid[96]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[97]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[113]_i_2_n_0 ),
        .I3(\valid[111]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [97]),
        .O(\valid[97]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[98]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[114]_i_2_n_0 ),
        .I3(\valid[111]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [98]),
        .O(\valid[98]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[99]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[115]_i_2_n_0 ),
        .I3(\valid[111]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [99]),
        .O(\valid[99]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \valid[9]_i_1 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\valid[121]_i_2_n_0 ),
        .I3(\valid[15]_i_2_n_0 ),
        .I4(\icache/state_reg_n_0_[2] ),
        .I5(\icache/valid [9]),
        .O(\valid[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_adr_out[0]_INST_0 
       (.I0(\dmem_if_outputs[adr] [0]),
        .I1(\arbiter/state [1]),
        .O(wb_adr_out[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_adr_out[1]_INST_0 
       (.I0(\dmem_if_outputs[adr] [1]),
        .I1(\arbiter/state [1]),
        .O(wb_adr_out[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[0]_INST_0 
       (.I0(\dmem_if_outputs[dat] [0]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[10]_INST_0 
       (.I0(\dmem_if_outputs[dat] [10]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[11]_INST_0 
       (.I0(\dmem_if_outputs[dat] [11]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[12]_INST_0 
       (.I0(\dmem_if_outputs[dat] [12]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[13]_INST_0 
       (.I0(\dmem_if_outputs[dat] [13]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[14]_INST_0 
       (.I0(\dmem_if_outputs[dat] [14]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[15]_INST_0 
       (.I0(\dmem_if_outputs[dat] [15]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[16]_INST_0 
       (.I0(\dmem_if_outputs[dat] [16]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[17]_INST_0 
       (.I0(\dmem_if_outputs[dat] [17]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[18]_INST_0 
       (.I0(\dmem_if_outputs[dat] [18]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[19]_INST_0 
       (.I0(\dmem_if_outputs[dat] [19]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[1]_INST_0 
       (.I0(\dmem_if_outputs[dat] [1]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[20]_INST_0 
       (.I0(\dmem_if_outputs[dat] [20]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[21]_INST_0 
       (.I0(\dmem_if_outputs[dat] [21]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[22]_INST_0 
       (.I0(\dmem_if_outputs[dat] [22]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[23]_INST_0 
       (.I0(\dmem_if_outputs[dat] [23]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[24]_INST_0 
       (.I0(\dmem_if_outputs[dat] [24]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[25]_INST_0 
       (.I0(\dmem_if_outputs[dat] [25]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[26]_INST_0 
       (.I0(\dmem_if_outputs[dat] [26]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[27]_INST_0 
       (.I0(\dmem_if_outputs[dat] [27]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[28]_INST_0 
       (.I0(\dmem_if_outputs[dat] [28]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[29]_INST_0 
       (.I0(\dmem_if_outputs[dat] [29]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[2]_INST_0 
       (.I0(\dmem_if_outputs[dat] [2]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[30]_INST_0 
       (.I0(\dmem_if_outputs[dat] [30]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[31]_INST_0 
       (.I0(\dmem_if_outputs[dat] [31]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[3]_INST_0 
       (.I0(\dmem_if_outputs[dat] [3]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[4]_INST_0 
       (.I0(\dmem_if_outputs[dat] [4]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[5]_INST_0 
       (.I0(\dmem_if_outputs[dat] [5]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[6]_INST_0 
       (.I0(\dmem_if_outputs[dat] [6]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[7]_INST_0 
       (.I0(\dmem_if_outputs[dat] [7]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[8]_INST_0 
       (.I0(\dmem_if_outputs[dat] [8]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_dat_out[9]_INST_0 
       (.I0(\dmem_if_outputs[dat] [9]),
        .I1(\arbiter/state [1]),
        .O(wb_dat_out[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][0]_i_1 
       (.I0(dmem_address_p[0]),
        .I1(\processor/ex_rd_data [0]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair140" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \wb_outputs[adr][10]_i_1 
       (.I0(\icache/cl_load_address [10]),
        .I1(imem_address[10]),
        .I2(\icache/state_reg_n_0_[2] ),
        .O(wb_outputs));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][10]_i_1__0 
       (.I0(dmem_address_p[10]),
        .I1(\processor/ex_rd_data [10]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair140" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \wb_outputs[adr][11]_i_1 
       (.I0(\icache/cl_load_address [11]),
        .I1(imem_address[11]),
        .I2(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][11]_i_1__0 
       (.I0(dmem_address_p[11]),
        .I1(\processor/ex_rd_data [11]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][12]_i_1 
       (.I0(dmem_address_p[12]),
        .I1(\processor/ex_rd_data [12]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00ACAC)) 
    \wb_outputs[adr][12]_i_1__0 
       (.I0(pc[12]),
        .I1(pc_next[12]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/cl_load_address [12]),
        .I4(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][12]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][13]_i_1 
       (.I0(dmem_address_p[13]),
        .I1(\processor/ex_rd_data [13]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00ACAC)) 
    \wb_outputs[adr][13]_i_1__0 
       (.I0(pc[13]),
        .I1(pc_next[13]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/cl_load_address [13]),
        .I4(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][13]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair135" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \wb_outputs[adr][14]_i_1 
       (.I0(\icache/cl_load_address [14]),
        .I1(imem_address[14]),
        .I2(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][14]_i_1__0 
       (.I0(dmem_address_p[14]),
        .I1(\processor/ex_rd_data [14]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][15]_i_1 
       (.I0(dmem_address_p[15]),
        .I1(\processor/ex_rd_data [15]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00ACAC)) 
    \wb_outputs[adr][15]_i_1__0 
       (.I0(pc[15]),
        .I1(pc_next[15]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/cl_load_address [15]),
        .I4(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][15]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][16]_i_1 
       (.I0(dmem_address_p[16]),
        .I1(\processor/ex_rd_data [16]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00ACAC)) 
    \wb_outputs[adr][16]_i_1__0 
       (.I0(pc[16]),
        .I1(pc_next[16]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/cl_load_address [16]),
        .I4(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][16]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair135" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \wb_outputs[adr][17]_i_1 
       (.I0(\icache/cl_load_address [17]),
        .I1(imem_address[17]),
        .I2(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][17]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][17]_i_1__0 
       (.I0(dmem_address_p[17]),
        .I1(\processor/ex_rd_data [17]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][18]_i_1 
       (.I0(dmem_address_p[18]),
        .I1(\processor/ex_rd_data [18]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00ACAC)) 
    \wb_outputs[adr][18]_i_1__0 
       (.I0(pc[18]),
        .I1(pc_next[18]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/cl_load_address [18]),
        .I4(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][18]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][19]_i_1 
       (.I0(dmem_address_p[19]),
        .I1(\processor/ex_rd_data [19]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00ACAC)) 
    \wb_outputs[adr][19]_i_1__0 
       (.I0(pc[19]),
        .I1(pc_next[19]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/cl_load_address [19]),
        .I4(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][19]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][1]_i_1 
       (.I0(dmem_address_p[1]),
        .I1(\processor/ex_rd_data [1]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair101" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \wb_outputs[adr][20]_i_1 
       (.I0(\icache/cl_load_address [20]),
        .I1(imem_address[20]),
        .I2(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][20]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][20]_i_1__0 
       (.I0(dmem_address_p[20]),
        .I1(\processor/ex_rd_data [20]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][21]_i_1 
       (.I0(dmem_address_p[21]),
        .I1(\processor/ex_rd_data [21]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00ACAC)) 
    \wb_outputs[adr][21]_i_1__0 
       (.I0(pc[21]),
        .I1(pc_next[21]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/cl_load_address [21]),
        .I4(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][21]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][22]_i_1 
       (.I0(dmem_address_p[22]),
        .I1(\processor/ex_rd_data [22]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00ACAC)) 
    \wb_outputs[adr][22]_i_1__0 
       (.I0(pc[22]),
        .I1(pc_next[22]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/cl_load_address [22]),
        .I4(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][22]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair101" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \wb_outputs[adr][23]_i_1 
       (.I0(\icache/cl_load_address [23]),
        .I1(imem_address[23]),
        .I2(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][23]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][23]_i_1__0 
       (.I0(dmem_address_p[23]),
        .I1(\processor/ex_rd_data [23]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][24]_i_1 
       (.I0(dmem_address_p[24]),
        .I1(\processor/ex_rd_data [24]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00ACAC)) 
    \wb_outputs[adr][24]_i_1__0 
       (.I0(pc[24]),
        .I1(pc_next[24]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/cl_load_address [24]),
        .I4(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][24]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][25]_i_1 
       (.I0(dmem_address_p[25]),
        .I1(\processor/ex_rd_data [25]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00ACAC)) 
    \wb_outputs[adr][25]_i_1__0 
       (.I0(pc[25]),
        .I1(pc_next[25]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/cl_load_address [25]),
        .I4(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][25]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair94" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \wb_outputs[adr][26]_i_1 
       (.I0(\icache/cl_load_address [26]),
        .I1(imem_address[26]),
        .I2(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][26]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][26]_i_1__0 
       (.I0(dmem_address_p[26]),
        .I1(\processor/ex_rd_data [26]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][27]_i_1 
       (.I0(dmem_address_p[27]),
        .I1(\processor/ex_rd_data [27]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00ACAC)) 
    \wb_outputs[adr][27]_i_1__0 
       (.I0(pc[27]),
        .I1(pc_next[27]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/cl_load_address [27]),
        .I4(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][27]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][28]_i_1 
       (.I0(dmem_address_p[28]),
        .I1(\processor/ex_rd_data [28]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00ACAC)) 
    \wb_outputs[adr][28]_i_1__0 
       (.I0(pc[28]),
        .I1(pc_next[28]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/cl_load_address [28]),
        .I4(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][28]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair94" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \wb_outputs[adr][29]_i_1 
       (.I0(\icache/cl_load_address [29]),
        .I1(imem_address[29]),
        .I2(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][29]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][29]_i_1__0 
       (.I0(dmem_address_p[29]),
        .I1(\processor/ex_rd_data [29]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][2]_i_1 
       (.I0(dmem_address_p[2]),
        .I1(\processor/ex_rd_data [2]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair195" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_outputs[adr][2]_i_1__0 
       (.I0(\icache/state_reg_n_0_[2] ),
        .I1(\icache/cl_current_word_reg_n_0_ ),
        .O(\wb_outputs[adr][2]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][30]_i_1 
       (.I0(dmem_address_p[30]),
        .I1(\processor/ex_rd_data [30]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00ACAC)) 
    \wb_outputs[adr][30]_i_1__0 
       (.I0(pc[30]),
        .I1(pc_next[30]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/cl_load_address [30]),
        .I4(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][30]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    \wb_outputs[adr][31]_i_1 
       (.I0(\dmem_if/state_reg_n_0_[1] ),
        .I1(\dmem_if/state_reg_n_0_ ),
        .I2(\wb_outputs[adr][31]_i_3_n_0 ),
        .I3(reset),
        .O(\wb_outputs[adr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00001011)) 
    \wb_outputs[adr][31]_i_1__0 
       (.I0(\icache/state_reg_n_0_[1] ),
        .I1(\icache/state_reg_n_0_ ),
        .I2(\icache/state_reg_n_0_[2] ),
        .I3(\icache/cache_hit ),
        .I4(reset),
        .O(\wb_outputs[adr][31]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][31]_i_2 
       (.I0(dmem_address_p[31]),
        .I1(\processor/ex_rd_data [31]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00ACAC)) 
    \wb_outputs[adr][31]_i_2__0 
       (.I0(pc[31]),
        .I1(pc_next[31]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/cl_load_address [31]),
        .I4(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][31]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAABAFFFFAABAAAAA)) 
    \wb_outputs[adr][31]_i_3 
       (.I0(dmem_write_req),
        .I1(\mem_op[2]_i_5_n_0 ),
        .I2(\processor/ex_mem_op [1]),
        .I3(\processor/ex_mem_op [2]),
        .I4(\processor/memory/p_1_in ),
        .I5(\processor/dmem_read_req_p ),
        .O(\wb_outputs[adr][31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][3]_i_1 
       (.I0(dmem_address_p[3]),
        .I1(\processor/ex_rd_data [3]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair195" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \wb_outputs[adr][3]_i_1__0 
       (.I0(\icache/state_reg_n_0_[2] ),
        .I1(\icache/cl_current_word_reg_n_0_[1] ),
        .O(\wb_outputs[adr][3]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair145" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \wb_outputs[adr][4]_i_1 
       (.I0(\icache/cl_load_address [4]),
        .I1(imem_address[4]),
        .I2(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][4]_i_1__0 
       (.I0(dmem_address_p[4]),
        .I1(\processor/ex_rd_data [4]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair145" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \wb_outputs[adr][5]_i_1 
       (.I0(\icache/cl_load_address [5]),
        .I1(imem_address[5]),
        .I2(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][5]_i_1__0 
       (.I0(dmem_address_p[5]),
        .I1(\processor/ex_rd_data [5]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][6]_i_1 
       (.I0(dmem_address_p[6]),
        .I1(\processor/ex_rd_data [6]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00ACAC)) 
    \wb_outputs[adr][6]_i_1__0 
       (.I0(pc[6]),
        .I1(pc_next[6]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/cl_load_address [6]),
        .I4(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][6]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][7]_i_1 
       (.I0(dmem_address_p[7]),
        .I1(\processor/ex_rd_data [7]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00ACAC)) 
    \wb_outputs[adr][7]_i_1__0 
       (.I0(pc[7]),
        .I1(pc_next[7]),
        .I2(\processor/fetch/cancel_fetch ),
        .I3(\icache/cl_load_address [7]),
        .I4(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][7]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \wb_outputs[adr][8]_i_1 
       (.I0(\icache/cl_load_address [8]),
        .I1(imem_address[8]),
        .I2(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][8]_i_1__0 
       (.I0(dmem_address_p[8]),
        .I1(\processor/ex_rd_data [8]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \wb_outputs[adr][9]_i_1 
       (.I0(\icache/cl_load_address [9]),
        .I1(imem_address[9]),
        .I2(\icache/state_reg_n_0_[2] ),
        .O(\wb_outputs[adr][9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0CAA)) 
    \wb_outputs[adr][9]_i_1__0 
       (.I0(dmem_address_p[9]),
        .I1(\processor/ex_rd_data [9]),
        .I2(\dmem_address_p[31]_i_2_n_0 ),
        .I3(\processor/memory/p_1_in ),
        .O(dmem_address__0[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h37370500)) 
    \wb_outputs[cyc]_i_1 
       (.I0(\dmem_if/state_reg_n_0_[1] ),
        .I1(dmem_if_inputs),
        .I2(\dmem_if/state_reg_n_0_ ),
        .I3(\wb_outputs[adr][31]_i_3_n_0 ),
        .I4(dmem_if_outputs),
        .O(\wb_outputs[cyc]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0F110FFF00110000)) 
    \wb_outputs[cyc]_i_1__0 
       (.I0(\icache/state_reg_n_0_[1] ),
        .I1(\icache/cache_hit ),
        .I2(\wb_outputs[cyc]_i_2_n_0 ),
        .I3(\icache/state_reg_n_0_[2] ),
        .I4(\wb_outputs[cyc]_i_3_n_0 ),
        .I5(icache_outputs),
        .O(\wb_outputs[cyc]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h20000000)) 
    \wb_outputs[cyc]_i_2 
       (.I0(\icache/state_reg_n_0_ ),
        .I1(\icache/cl_current_word_reg_n_0_[2] ),
        .I2(\icache/cl_current_word_reg_n_0_ ),
        .I3(\icache/cl_current_word_reg_n_0_[1] ),
        .I4(icache_inputs),
        .O(\wb_outputs[cyc]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h40004000400040FF)) 
    \wb_outputs[cyc]_i_3 
       (.I0(\arbiter/state [1]),
        .I1(\arbiter/state [0]),
        .I2(wb_ack_in),
        .I3(\icache/state_reg_n_0_[1] ),
        .I4(\icache/state_reg_n_0_ ),
        .I5(\icache/cache_hit ),
        .O(\wb_outputs[cyc]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00D8)) 
    \wb_outputs[dat][0]_i_1 
       (.I0(\processor/memory/p_1_in ),
        .I1(\processor/ex_dmem_data_out [0]),
        .I2(dmem_data_out_p[0]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .O(\wb_outputs[dat][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000D8FFD800)) 
    \wb_outputs[dat][10]_i_1 
       (.I0(\processor/memory/p_1_in ),
        .I1(\processor/ex_dmem_data_out [2]),
        .I2(dmem_data_out_p[2]),
        .I3(\dmem_data_out[23]_i_3_n_0 ),
        .I4(dmem_data_in[10]),
        .I5(\dmem_data_out[23]_i_4_n_0 ),
        .O(SHIFT_LEFT[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \wb_outputs[dat][10]_i_2 
       (.I0(dmem_data_out_p[10]),
        .I1(\processor/ex_dmem_data_out [10]),
        .I2(\processor/memory/p_1_in ),
        .O(dmem_data_in[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000D8FFD800)) 
    \wb_outputs[dat][11]_i_1 
       (.I0(\processor/memory/p_1_in ),
        .I1(\processor/ex_dmem_data_out [3]),
        .I2(dmem_data_out_p[3]),
        .I3(\dmem_data_out[23]_i_3_n_0 ),
        .I4(dmem_data_in[11]),
        .I5(\dmem_data_out[23]_i_4_n_0 ),
        .O(SHIFT_LEFT[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \wb_outputs[dat][11]_i_2 
       (.I0(dmem_data_out_p[11]),
        .I1(\processor/ex_dmem_data_out [11]),
        .I2(\processor/memory/p_1_in ),
        .O(dmem_data_in[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000D8FFD800)) 
    \wb_outputs[dat][12]_i_1 
       (.I0(\processor/memory/p_1_in ),
        .I1(\processor/ex_dmem_data_out [4]),
        .I2(dmem_data_out_p[4]),
        .I3(\dmem_data_out[23]_i_3_n_0 ),
        .I4(dmem_data_in[12]),
        .I5(\dmem_data_out[23]_i_4_n_0 ),
        .O(SHIFT_LEFT[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \wb_outputs[dat][12]_i_2 
       (.I0(dmem_data_out_p[12]),
        .I1(\processor/ex_dmem_data_out [12]),
        .I2(\processor/memory/p_1_in ),
        .O(dmem_data_in[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000D8FFD800)) 
    \wb_outputs[dat][13]_i_1 
       (.I0(\processor/memory/p_1_in ),
        .I1(\processor/ex_dmem_data_out [5]),
        .I2(dmem_data_out_p[5]),
        .I3(\dmem_data_out[23]_i_3_n_0 ),
        .I4(dmem_data_in[13]),
        .I5(\dmem_data_out[23]_i_4_n_0 ),
        .O(SHIFT_LEFT[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \wb_outputs[dat][13]_i_2 
       (.I0(dmem_data_out_p[13]),
        .I1(\processor/ex_dmem_data_out [13]),
        .I2(\processor/memory/p_1_in ),
        .O(dmem_data_in[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000D8FFD800)) 
    \wb_outputs[dat][14]_i_1 
       (.I0(\processor/memory/p_1_in ),
        .I1(\processor/ex_dmem_data_out [6]),
        .I2(dmem_data_out_p[6]),
        .I3(\dmem_data_out[23]_i_3_n_0 ),
        .I4(dmem_data_in[14]),
        .I5(\dmem_data_out[23]_i_4_n_0 ),
        .O(SHIFT_LEFT[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \wb_outputs[dat][14]_i_2 
       (.I0(dmem_data_out_p[14]),
        .I1(\processor/ex_dmem_data_out [14]),
        .I2(\processor/memory/p_1_in ),
        .O(dmem_data_in[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000D8FFD800)) 
    \wb_outputs[dat][15]_i_1 
       (.I0(\processor/memory/p_1_in ),
        .I1(\processor/ex_dmem_data_out [7]),
        .I2(dmem_data_out_p[7]),
        .I3(\dmem_data_out[23]_i_3_n_0 ),
        .I4(dmem_data_in[15]),
        .I5(\dmem_data_out[23]_i_4_n_0 ),
        .O(SHIFT_LEFT[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \wb_outputs[dat][15]_i_2 
       (.I0(dmem_data_out_p[15]),
        .I1(\processor/ex_dmem_data_out [15]),
        .I2(\processor/memory/p_1_in ),
        .O(dmem_data_in[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00D8FFFF00D80000)) 
    \wb_outputs[dat][16]_i_1 
       (.I0(\processor/memory/p_1_in ),
        .I1(\processor/ex_dmem_data_out [8]),
        .I2(dmem_data_out_p[8]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .I4(\dmem_data_out[23]_i_3_n_0 ),
        .I5(\wb_outputs[dat][24]_i_2_n_0 ),
        .O(SHIFT_LEFT[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00D8FFFF00D80000)) 
    \wb_outputs[dat][17]_i_1 
       (.I0(\processor/memory/p_1_in ),
        .I1(\processor/ex_dmem_data_out [9]),
        .I2(dmem_data_out_p[9]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .I4(\dmem_data_out[23]_i_3_n_0 ),
        .I5(\wb_outputs[dat][25]_i_2_n_0 ),
        .O(SHIFT_LEFT[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00D8FFFF00D80000)) 
    \wb_outputs[dat][18]_i_1 
       (.I0(\processor/memory/p_1_in ),
        .I1(\processor/ex_dmem_data_out [10]),
        .I2(dmem_data_out_p[10]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .I4(\dmem_data_out[23]_i_3_n_0 ),
        .I5(\wb_outputs[dat][26]_i_2_n_0 ),
        .O(SHIFT_LEFT[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00D8FFFF00D80000)) 
    \wb_outputs[dat][19]_i_1 
       (.I0(\processor/memory/p_1_in ),
        .I1(\processor/ex_dmem_data_out [11]),
        .I2(dmem_data_out_p[11]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .I4(\dmem_data_out[23]_i_3_n_0 ),
        .I5(\wb_outputs[dat][27]_i_2_n_0 ),
        .O(SHIFT_LEFT[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00D8)) 
    \wb_outputs[dat][1]_i_1 
       (.I0(\processor/memory/p_1_in ),
        .I1(\processor/ex_dmem_data_out [1]),
        .I2(dmem_data_out_p[1]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .O(\wb_outputs[dat][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00D8FFFF00D80000)) 
    \wb_outputs[dat][20]_i_1 
       (.I0(\processor/memory/p_1_in ),
        .I1(\processor/ex_dmem_data_out [12]),
        .I2(dmem_data_out_p[12]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .I4(\dmem_data_out[23]_i_3_n_0 ),
        .I5(\wb_outputs[dat][28]_i_2_n_0 ),
        .O(SHIFT_LEFT[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00D8FFFF00D80000)) 
    \wb_outputs[dat][21]_i_1 
       (.I0(\processor/memory/p_1_in ),
        .I1(\processor/ex_dmem_data_out [13]),
        .I2(dmem_data_out_p[13]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .I4(\dmem_data_out[23]_i_3_n_0 ),
        .I5(\wb_outputs[dat][29]_i_2_n_0 ),
        .O(SHIFT_LEFT[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00D8FFFF00D80000)) 
    \wb_outputs[dat][22]_i_1 
       (.I0(\processor/memory/p_1_in ),
        .I1(\processor/ex_dmem_data_out [14]),
        .I2(dmem_data_out_p[14]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .I4(\dmem_data_out[23]_i_3_n_0 ),
        .I5(\wb_outputs[dat][30]_i_2_n_0 ),
        .O(SHIFT_LEFT[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00D8FFFF00D80000)) 
    \wb_outputs[dat][23]_i_1 
       (.I0(\processor/memory/p_1_in ),
        .I1(\processor/ex_dmem_data_out [15]),
        .I2(dmem_data_out_p[15]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .I4(\dmem_data_out[23]_i_3_n_0 ),
        .I5(\wb_outputs[dat][31]_i_3_n_0 ),
        .O(SHIFT_LEFT[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair170" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \wb_outputs[dat][24]_i_1 
       (.I0(\wb_outputs[dat][24]_i_2_n_0 ),
        .I1(\dmem_data_out[23]_i_3_n_0 ),
        .I2(\wb_outputs[dat][24]_i_3_n_0 ),
        .O(SHIFT_LEFT[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFCFC0C0AFA0AFA0)) 
    \wb_outputs[dat][24]_i_2 
       (.I0(dmem_data_out_p[0]),
        .I1(\processor/ex_dmem_data_out [0]),
        .I2(\dmem_data_out[23]_i_4_n_0 ),
        .I3(dmem_data_out_p[16]),
        .I4(\processor/ex_dmem_data_out [16]),
        .I5(\processor/memory/p_1_in ),
        .O(\wb_outputs[dat][24]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFCFC0C0AFA0AFA0)) 
    \wb_outputs[dat][24]_i_3 
       (.I0(dmem_data_out_p[8]),
        .I1(\processor/ex_dmem_data_out [8]),
        .I2(\dmem_data_out[23]_i_4_n_0 ),
        .I3(dmem_data_out_p[24]),
        .I4(\processor/ex_dmem_data_out [24]),
        .I5(\processor/memory/p_1_in ),
        .O(\wb_outputs[dat][24]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair170" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \wb_outputs[dat][25]_i_1 
       (.I0(\wb_outputs[dat][25]_i_2_n_0 ),
        .I1(\dmem_data_out[23]_i_3_n_0 ),
        .I2(\wb_outputs[dat][25]_i_3_n_0 ),
        .O(SHIFT_LEFT[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFCFC0C0AFA0AFA0)) 
    \wb_outputs[dat][25]_i_2 
       (.I0(dmem_data_out_p[1]),
        .I1(\processor/ex_dmem_data_out [1]),
        .I2(\dmem_data_out[23]_i_4_n_0 ),
        .I3(dmem_data_out_p[17]),
        .I4(\processor/ex_dmem_data_out [17]),
        .I5(\processor/memory/p_1_in ),
        .O(\wb_outputs[dat][25]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFCFC0C0AFA0AFA0)) 
    \wb_outputs[dat][25]_i_3 
       (.I0(dmem_data_out_p[9]),
        .I1(\processor/ex_dmem_data_out [9]),
        .I2(\dmem_data_out[23]_i_4_n_0 ),
        .I3(dmem_data_out_p[25]),
        .I4(\processor/ex_dmem_data_out [25]),
        .I5(\processor/memory/p_1_in ),
        .O(\wb_outputs[dat][25]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair157" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \wb_outputs[dat][26]_i_1 
       (.I0(\wb_outputs[dat][26]_i_2_n_0 ),
        .I1(\dmem_data_out[23]_i_3_n_0 ),
        .I2(\wb_outputs[dat][26]_i_3_n_0 ),
        .O(SHIFT_LEFT[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFCFC0C0AFA0AFA0)) 
    \wb_outputs[dat][26]_i_2 
       (.I0(dmem_data_out_p[2]),
        .I1(\processor/ex_dmem_data_out [2]),
        .I2(\dmem_data_out[23]_i_4_n_0 ),
        .I3(dmem_data_out_p[18]),
        .I4(\processor/ex_dmem_data_out [18]),
        .I5(\processor/memory/p_1_in ),
        .O(\wb_outputs[dat][26]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFCFC0C0AFA0AFA0)) 
    \wb_outputs[dat][26]_i_3 
       (.I0(dmem_data_out_p[10]),
        .I1(\processor/ex_dmem_data_out [10]),
        .I2(\dmem_data_out[23]_i_4_n_0 ),
        .I3(dmem_data_out_p[26]),
        .I4(\processor/ex_dmem_data_out [26]),
        .I5(\processor/memory/p_1_in ),
        .O(\wb_outputs[dat][26]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair157" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \wb_outputs[dat][27]_i_1 
       (.I0(\wb_outputs[dat][27]_i_2_n_0 ),
        .I1(\dmem_data_out[23]_i_3_n_0 ),
        .I2(\wb_outputs[dat][27]_i_3_n_0 ),
        .O(SHIFT_LEFT[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFCFC0C0AFA0AFA0)) 
    \wb_outputs[dat][27]_i_2 
       (.I0(dmem_data_out_p[3]),
        .I1(\processor/ex_dmem_data_out [3]),
        .I2(\dmem_data_out[23]_i_4_n_0 ),
        .I3(dmem_data_out_p[19]),
        .I4(\processor/ex_dmem_data_out [19]),
        .I5(\processor/memory/p_1_in ),
        .O(\wb_outputs[dat][27]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFCFC0C0AFA0AFA0)) 
    \wb_outputs[dat][27]_i_3 
       (.I0(dmem_data_out_p[11]),
        .I1(\processor/ex_dmem_data_out [11]),
        .I2(\dmem_data_out[23]_i_4_n_0 ),
        .I3(dmem_data_out_p[27]),
        .I4(\processor/ex_dmem_data_out [27]),
        .I5(\processor/memory/p_1_in ),
        .O(\wb_outputs[dat][27]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair156" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \wb_outputs[dat][28]_i_1 
       (.I0(\wb_outputs[dat][28]_i_2_n_0 ),
        .I1(\dmem_data_out[23]_i_3_n_0 ),
        .I2(\wb_outputs[dat][28]_i_3_n_0 ),
        .O(SHIFT_LEFT[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFCFC0C0AFA0AFA0)) 
    \wb_outputs[dat][28]_i_2 
       (.I0(dmem_data_out_p[4]),
        .I1(\processor/ex_dmem_data_out [4]),
        .I2(\dmem_data_out[23]_i_4_n_0 ),
        .I3(dmem_data_out_p[20]),
        .I4(\processor/ex_dmem_data_out [20]),
        .I5(\processor/memory/p_1_in ),
        .O(\wb_outputs[dat][28]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFCFC0C0AFA0AFA0)) 
    \wb_outputs[dat][28]_i_3 
       (.I0(dmem_data_out_p[12]),
        .I1(\processor/ex_dmem_data_out [12]),
        .I2(\dmem_data_out[23]_i_4_n_0 ),
        .I3(dmem_data_out_p[28]),
        .I4(\processor/ex_dmem_data_out [28]),
        .I5(\processor/memory/p_1_in ),
        .O(\wb_outputs[dat][28]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair156" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \wb_outputs[dat][29]_i_1 
       (.I0(\wb_outputs[dat][29]_i_2_n_0 ),
        .I1(\dmem_data_out[23]_i_3_n_0 ),
        .I2(\wb_outputs[dat][29]_i_3_n_0 ),
        .O(SHIFT_LEFT[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFCFC0C0AFA0AFA0)) 
    \wb_outputs[dat][29]_i_2 
       (.I0(dmem_data_out_p[5]),
        .I1(\processor/ex_dmem_data_out [5]),
        .I2(\dmem_data_out[23]_i_4_n_0 ),
        .I3(dmem_data_out_p[21]),
        .I4(\processor/ex_dmem_data_out [21]),
        .I5(\processor/memory/p_1_in ),
        .O(\wb_outputs[dat][29]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFCFC0C0AFA0AFA0)) 
    \wb_outputs[dat][29]_i_3 
       (.I0(dmem_data_out_p[13]),
        .I1(\processor/ex_dmem_data_out [13]),
        .I2(\dmem_data_out[23]_i_4_n_0 ),
        .I3(dmem_data_out_p[29]),
        .I4(\processor/ex_dmem_data_out [29]),
        .I5(\processor/memory/p_1_in ),
        .O(\wb_outputs[dat][29]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00D8)) 
    \wb_outputs[dat][2]_i_1 
       (.I0(\processor/memory/p_1_in ),
        .I1(\processor/ex_dmem_data_out [2]),
        .I2(dmem_data_out_p[2]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .O(\wb_outputs[dat][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair155" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \wb_outputs[dat][30]_i_1 
       (.I0(\wb_outputs[dat][30]_i_2_n_0 ),
        .I1(\dmem_data_out[23]_i_3_n_0 ),
        .I2(\wb_outputs[dat][30]_i_3_n_0 ),
        .O(SHIFT_LEFT[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFCFC0C0AFA0AFA0)) 
    \wb_outputs[dat][30]_i_2 
       (.I0(dmem_data_out_p[6]),
        .I1(\processor/ex_dmem_data_out [6]),
        .I2(\dmem_data_out[23]_i_4_n_0 ),
        .I3(dmem_data_out_p[22]),
        .I4(\processor/ex_dmem_data_out [22]),
        .I5(\processor/memory/p_1_in ),
        .O(\wb_outputs[dat][30]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFCFC0C0AFA0AFA0)) 
    \wb_outputs[dat][30]_i_3 
       (.I0(dmem_data_out_p[14]),
        .I1(\processor/ex_dmem_data_out [14]),
        .I2(\dmem_data_out[23]_i_4_n_0 ),
        .I3(dmem_data_out_p[30]),
        .I4(\processor/ex_dmem_data_out [30]),
        .I5(\processor/memory/p_1_in ),
        .O(\wb_outputs[dat][30]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    \wb_outputs[dat][31]_i_1 
       (.I0(\dmem_if/state_reg_n_0_[1] ),
        .I1(\dmem_if/state_reg_n_0_ ),
        .I2(dmem_write_req),
        .I3(reset),
        .O(\wb_outputs[dat][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair155" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \wb_outputs[dat][31]_i_2 
       (.I0(\wb_outputs[dat][31]_i_3_n_0 ),
        .I1(\dmem_data_out[23]_i_3_n_0 ),
        .I2(\wb_outputs[dat][31]_i_4_n_0 ),
        .O(SHIFT_LEFT[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFCFC0C0AFA0AFA0)) 
    \wb_outputs[dat][31]_i_3 
       (.I0(dmem_data_out_p[7]),
        .I1(\processor/ex_dmem_data_out [7]),
        .I2(\dmem_data_out[23]_i_4_n_0 ),
        .I3(dmem_data_out_p[23]),
        .I4(\processor/ex_dmem_data_out [23]),
        .I5(\processor/memory/p_1_in ),
        .O(\wb_outputs[dat][31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFCFC0C0AFA0AFA0)) 
    \wb_outputs[dat][31]_i_4 
       (.I0(dmem_data_out_p[15]),
        .I1(\processor/ex_dmem_data_out [15]),
        .I2(\dmem_data_out[23]_i_4_n_0 ),
        .I3(dmem_data_out_p[31]),
        .I4(\processor/ex_dmem_data_out [31]),
        .I5(\processor/memory/p_1_in ),
        .O(\wb_outputs[dat][31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00D8)) 
    \wb_outputs[dat][3]_i_1 
       (.I0(\processor/memory/p_1_in ),
        .I1(\processor/ex_dmem_data_out [3]),
        .I2(dmem_data_out_p[3]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .O(\wb_outputs[dat][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00D8)) 
    \wb_outputs[dat][4]_i_1 
       (.I0(\processor/memory/p_1_in ),
        .I1(\processor/ex_dmem_data_out [4]),
        .I2(dmem_data_out_p[4]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .O(\wb_outputs[dat][4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00D8)) 
    \wb_outputs[dat][5]_i_1 
       (.I0(\processor/memory/p_1_in ),
        .I1(\processor/ex_dmem_data_out [5]),
        .I2(dmem_data_out_p[5]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .O(\wb_outputs[dat][5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00D8)) 
    \wb_outputs[dat][6]_i_1 
       (.I0(\processor/memory/p_1_in ),
        .I1(\processor/ex_dmem_data_out [6]),
        .I2(dmem_data_out_p[6]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .O(\wb_outputs[dat][6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00100000)) 
    \wb_outputs[dat][7]_i_1 
       (.I0(\dmem_if/state_reg_n_0_[1] ),
        .I1(\dmem_if/state_reg_n_0_ ),
        .I2(dmem_write_req),
        .I3(reset),
        .I4(\dmem_data_out[23]_i_3_n_0 ),
        .O(\wb_outputs[dat][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00D8)) 
    \wb_outputs[dat][7]_i_2 
       (.I0(\processor/memory/p_1_in ),
        .I1(\processor/ex_dmem_data_out [7]),
        .I2(dmem_data_out_p[7]),
        .I3(\dmem_data_out[23]_i_4_n_0 ),
        .O(\wb_outputs[dat][7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000D8FFD800)) 
    \wb_outputs[dat][8]_i_1 
       (.I0(\processor/memory/p_1_in ),
        .I1(\processor/ex_dmem_data_out [0]),
        .I2(dmem_data_out_p[0]),
        .I3(\dmem_data_out[23]_i_3_n_0 ),
        .I4(dmem_data_in[8]),
        .I5(\dmem_data_out[23]_i_4_n_0 ),
        .O(SHIFT_LEFT[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \wb_outputs[dat][8]_i_2 
       (.I0(dmem_data_out_p[8]),
        .I1(\processor/ex_dmem_data_out [8]),
        .I2(\processor/memory/p_1_in ),
        .O(dmem_data_in[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000D8FFD800)) 
    \wb_outputs[dat][9]_i_1 
       (.I0(\processor/memory/p_1_in ),
        .I1(\processor/ex_dmem_data_out [1]),
        .I2(dmem_data_out_p[1]),
        .I3(\dmem_data_out[23]_i_3_n_0 ),
        .I4(dmem_data_in[9]),
        .I5(\dmem_data_out[23]_i_4_n_0 ),
        .O(SHIFT_LEFT[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \wb_outputs[dat][9]_i_2 
       (.I0(dmem_data_out_p[9]),
        .I1(\processor/ex_dmem_data_out [9]),
        .I2(\processor/memory/p_1_in ),
        .O(dmem_data_in[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000007D557DFF)) 
    \wb_outputs[sel][0]_i_1 
       (.I0(dmem_address[0]),
        .I1(\processor/ex_mem_size ),
        .I2(\processor/ex_dmem_data_size [1]),
        .I3(\processor/memory/p_1_in ),
        .I4(\processor/dmem_data_size_p [0]),
        .I5(dmem_address[1]),
        .O(\wb_outputs[sel][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000BEAABEFF)) 
    \wb_outputs[sel][1]_i_1 
       (.I0(dmem_address[0]),
        .I1(\processor/ex_mem_size ),
        .I2(\processor/ex_dmem_data_size [1]),
        .I3(\processor/memory/p_1_in ),
        .I4(\processor/dmem_data_size_p [0]),
        .I5(dmem_address[1]),
        .O(\wb_outputs[sel][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7D557DFF00000000)) 
    \wb_outputs[sel][2]_i_1 
       (.I0(dmem_address[0]),
        .I1(\processor/ex_mem_size ),
        .I2(\processor/ex_dmem_data_size [1]),
        .I3(\processor/memory/p_1_in ),
        .I4(\processor/dmem_data_size_p [0]),
        .I5(dmem_address[1]),
        .O(\wb_outputs[sel][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \wb_outputs[sel][3]_i_1 
       (.I0(\icache/cache_hit ),
        .O(\icache/p_1_in10_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA8A20802)) 
    \wb_outputs[sel][3]_i_1__0 
       (.I0(\wb_outputs[adr][31]_i_1_n_0 ),
        .I1(\processor/dmem_data_size_p [1]),
        .I2(\processor/memory/p_1_in ),
        .I3(\processor/dmem_data_size_p [0]),
        .I4(\processor/ex_mem_size ),
        .O(\wb_outputs[sel][3]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBEAABEFF00000000)) 
    \wb_outputs[sel][3]_i_2 
       (.I0(dmem_address[0]),
        .I1(\processor/ex_mem_size ),
        .I2(\processor/ex_dmem_data_size [1]),
        .I3(\processor/memory/p_1_in ),
        .I4(\processor/dmem_data_size_p [0]),
        .I5(dmem_address[1]),
        .O(\wb_outputs[sel][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair38" *) 
  LUT5 #(
    .INIT(32'hDF770300)) 
    \wb_outputs[stb]_i_1 
       (.I0(icache_inputs),
        .I1(\icache/state_reg_n_0_[1] ),
        .I2(\icache/state_reg_n_0_ ),
        .I3(\icache/state_reg_n_0_[2] ),
        .I4(\icache_outputs[stb] ),
        .O(\wb_outputs[stb]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF2F0020)) 
    \wb_outputs[we]_i_1 
       (.I0(dmem_write_req),
        .I1(\dmem_if/state_reg_n_0_[1] ),
        .I2(\wb_outputs[we]_i_2_n_0 ),
        .I3(reset),
        .I4(\dmem_if_outputs[we] ),
        .O(\wb_outputs[we]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000002222E222)) 
    \wb_outputs[we]_i_2 
       (.I0(\wb_outputs[adr][31]_i_3_n_0 ),
        .I1(\dmem_if/state_reg_n_0_[1] ),
        .I2(\arbiter/state [1]),
        .I3(wb_ack_in),
        .I4(\arbiter/state [0]),
        .I5(\dmem_if/state_reg_n_0_ ),
        .O(\wb_outputs[we]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    wb_we_out_INST_0
       (.I0(\arbiter/state [1]),
        .I1(\dmem_if_outputs[we] ),
        .O(wb_we_out));
endmodule
