module des3_area
   (desOut,
    desIn,
    key1,
    key2,
    key3,
    decrypt,
    roundSel,
    backdoor,
    clk);
  output backdoor;
  output [63:0]desOut;
  input [63:0]desIn;
  input [55:0]key1;
  input [55:0]key2;
  input [55:0]key3;
  input decrypt;
  input [5:0]roundSel;
  input clk;

  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const0>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const1>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire FP_R_reg_n_0_;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[42] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[43] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[44] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[45] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[46] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[47] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[48] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[49] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[50] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[51] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[52] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[53] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[54] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[55] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[56] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[57] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[58] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[59] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[60] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[61] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[62] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[63] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FP_R_reg_n_0_[64] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]R;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire clk;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire decrypt;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:0]desIn;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:0]desOut;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \desOut[62]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \desOut[62]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \desOut[63]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \desOut[63]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_100__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_100__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_100_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_101__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_101__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_101__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_101_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_102__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_102__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_102__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_102_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_103__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_103__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_103_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_104__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_104__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_104_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_105__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_105__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_105_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_106__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_106_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_107__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_107_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_108__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_108_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_109__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_109_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_10__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_10__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_10__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_10__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_10__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_10__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_10__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_110__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_110_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_111__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_111_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_112__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_112_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_113_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_114_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_115_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_116_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_117_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_118_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_119_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_11__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_11__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_11__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_11__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_11__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_11__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_11__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_120_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_121_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_122_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_123_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_124_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_125_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_126_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_127_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_128_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_129_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_12__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_12__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_12__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_12__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_12__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_12__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_12__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_130_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_131_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_13__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_13__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_13__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_13__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_13__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_13__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_13__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_14__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_14__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_14__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_14__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_14__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_14__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_14__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_15__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_15__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_15__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_15__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_15__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_15__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_15__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_16__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_16__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_16__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_16__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_16__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_16__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_16__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_17__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_17__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_17__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_17__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_17__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_17__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_17__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_18__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_18__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_18__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_18__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_18__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_18__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_18__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_19__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_19__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_19__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_19__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_19__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_19__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_19__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_20__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_20__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_20__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_20__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_20__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_20__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_20__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_21__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_21__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_21__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_21__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_21__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_21__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_21__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_22__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_22__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_22__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_22__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_22__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_22__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_22__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_23__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_23__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_23__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_23__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_23__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_23__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_23__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_24__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_24__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_24__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_24__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_24__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_24__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_24__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_24_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_25__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_25__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_25__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_25__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_25__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_25__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_25__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_25_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_26__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_26__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_26__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_26__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_26__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_26__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_26__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_26_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_27__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_27__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_27__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_27__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_27__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_27__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_27__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_27_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_28__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_28__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_28__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_28__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_28__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_28__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_28__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_28_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_29__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_29__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_29__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_29__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_29__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_29__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_29__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_29_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_30__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_30__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_30__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_30__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_30__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_30__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_30__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_30_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_31__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_31__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_31__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_31__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_31__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_31__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_31__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_31_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_32__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_32__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_32__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_32__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_32__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_32__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_32__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_32_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_33__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_33__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_33__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_33__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_33__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_33__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_33__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_33_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_34__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_34__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_34__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_34__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_34__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_34__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_34__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_34_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_35__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_35__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_35__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_35__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_35__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_35__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_35__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_35_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_36__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_36__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_36__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_36__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_36__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_36__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_36__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_36_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_37__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_37__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_37__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_37__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_37__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_37__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_37__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_37_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_38__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_38__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_38__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_38__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_38__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_38__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_38__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_38_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_39__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_39__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_39__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_39__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_39__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_39__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_39__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_39_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_40__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_40__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_40__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_40__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_40__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_40__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_40__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_40_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_41__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_41__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_41__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_41__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_41__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_41__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_41__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_41_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_42__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_42__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_42__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_42__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_42__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_42__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_42__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_42_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_43__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_43__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_43__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_43__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_43__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_43__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_43__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_43_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_44__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_44__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_44__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_44__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_44__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_44__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_44__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_44_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_45__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_45__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_45__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_45__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_45__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_45__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_45__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_45_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_46__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_46__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_46__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_46__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_46__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_46__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_46__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_46_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_47__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_47__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_47__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_47__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_47__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_47__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_47__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_47_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_48__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_48__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_48__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_48__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_48__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_48__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_48__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_48_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_49__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_49__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_49__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_49__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_49__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_49__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_49__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_49_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_50__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_50__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_50__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_50__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_50__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_50__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_50__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_50_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_51__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_51__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_51__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_51__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_51__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_51__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_51__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_51_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_52__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_52__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_52__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_52__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_52__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_52__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_52__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_52_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_53__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_53__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_53__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_53__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_53__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_53__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_53__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_53_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_54__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_54__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_54__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_54__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_54__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_54__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_54__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_54_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_55__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_55__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_55__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_55__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_55__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_55__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_55__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_55_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_56__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_56__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_56__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_56__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_56__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_56__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_56__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_56_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_57__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_57__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_57__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_57__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_57__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_57__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_57__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_57_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_58__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_58__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_58__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_58__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_58__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_58__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_58__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_58_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_59__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_59__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_59__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_59__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_59__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_59__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_59__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_59_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_60__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_60__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_60__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_60__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_60__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_60__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_60__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_60_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_61__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_61__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_61__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_61__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_61__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_61__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_61__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_61_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_62__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_62__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_62__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_62__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_62__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_62__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_62__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_62_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_63__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_63__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_63__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_63__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_63__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_63__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_63__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_63_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_64__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_64__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_64__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_64__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_64__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_64__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_64__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_64_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_65__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_65__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_65__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_65__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_65__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_65_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_66__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_66__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_66__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_66__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_66__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_66__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_66_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_67__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_67__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_67__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_67__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_67__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_67__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_67__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_67_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_68__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_68__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_68__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_68__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_68__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_68__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_68_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_69__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_69__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_69__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_69__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_69__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_69__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_69_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_70__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_70__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_70__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_70__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_70__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_70__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_70_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_71__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_71__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_71__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_71__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_71__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_71__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_71__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_71_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_72__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_72__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_72__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_72__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_72__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_72__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_72__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_72_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_73__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_73__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_73__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_73__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_73__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_73__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_73__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_73_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_74__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_74__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_74__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_74__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_74__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_74__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_74__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_74_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_75__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_75__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_75__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_75__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_75__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_75__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_75__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_75_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_76__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_76__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_76__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_76__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_76__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_76__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_76_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_77__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_77__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_77__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_77__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_77__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_77__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_77__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_77_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_78__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_78__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_78__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_78__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_78__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_78__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_78_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_79__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_79__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_79__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_79__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_79__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_79__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_79_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_7__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_7__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_7__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_7__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_7__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_7__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_7__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_80__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_80__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_80__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_80__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_80__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_80__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_80_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_81__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_81__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_81__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_81__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_81__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_81__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_81__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_81_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_82__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_82__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_82__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_82__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_82__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_82__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_82__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_82_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_83__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_83__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_83__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_83__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_83__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_83__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_83__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_83_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_84__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_84__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_84__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_84__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_84__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_84__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_84__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_84_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_85__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_85__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_85__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_85__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_85_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_86__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_86__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_86__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_86_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_87__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_87__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_87__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_87_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_88__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_88__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_88__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_88_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_89__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_89__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_89__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_89__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_89_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_8__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_8__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_8__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_8__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_8__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_8__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_8__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_90__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_90__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_90__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_90_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_91__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_91__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_91__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_91__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_91_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_92__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_92__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_92__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_92__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_92_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_93__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_93__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_93__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_93__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_93_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_94__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_94__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_94__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_94__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_94_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_95__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_95__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_95__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_95_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_96__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_96__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_96__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_96_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_97__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_97__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_97_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_98__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_98__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_98__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_98_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_99__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_99__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_99_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_9__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_9__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_9__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_9__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_9__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_9__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_9__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]key1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]key2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]key3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:0]roundSel;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u0/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/decrypt_int__2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/p_10_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/p_11_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/p_13_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/p_14_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/p_15_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/p_16_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/p_17_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/p_18_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/p_19_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/p_2_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/p_3_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/p_5_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/p_7_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/p_8_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/p_9_in ;

  assign backdoor =  \u1/p_9_in  ;

  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[7]),
        .Q(FP_R_reg_n_0_),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[15]),
        .Q(\FP_R_reg_n_0_[34] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[23]),
        .Q(\FP_R_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[31]),
        .Q(\FP_R_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[39]),
        .Q(\FP_R_reg_n_0_[37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[47]),
        .Q(\FP_R_reg_n_0_[38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[55]),
        .Q(\FP_R_reg_n_0_[39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[63]),
        .Q(\FP_R_reg_n_0_[40] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[5]),
        .Q(\FP_R_reg_n_0_[41] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[13]),
        .Q(\FP_R_reg_n_0_[42] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[21]),
        .Q(\FP_R_reg_n_0_[43] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[29]),
        .Q(\FP_R_reg_n_0_[44] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[37]),
        .Q(\FP_R_reg_n_0_[45] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[45]),
        .Q(\FP_R_reg_n_0_[46] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[53]),
        .Q(\FP_R_reg_n_0_[47] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[61]),
        .Q(\FP_R_reg_n_0_[48] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[3]),
        .Q(\FP_R_reg_n_0_[49] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[11]),
        .Q(\FP_R_reg_n_0_[50] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[19]),
        .Q(\FP_R_reg_n_0_[51] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[27]),
        .Q(\FP_R_reg_n_0_[52] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[35]),
        .Q(\FP_R_reg_n_0_[53] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[43]),
        .Q(\FP_R_reg_n_0_[54] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[51]),
        .Q(\FP_R_reg_n_0_[55] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[59]),
        .Q(\FP_R_reg_n_0_[56] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[1]),
        .Q(\FP_R_reg_n_0_[57] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[9]),
        .Q(\FP_R_reg_n_0_[58] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[17]),
        .Q(\FP_R_reg_n_0_[59] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[25]),
        .Q(\FP_R_reg_n_0_[60] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[33]),
        .Q(\FP_R_reg_n_0_[61] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[41]),
        .Q(\FP_R_reg_n_0_[62] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[49]),
        .Q(\FP_R_reg_n_0_[63] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \FP_R_reg[64] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[57]),
        .Q(\FP_R_reg_n_0_[64] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND
       (.G(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[12]),
        .Q(R[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[20]),
        .Q(R[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[28]),
        .Q(R[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[36]),
        .Q(R[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[44]),
        .Q(R[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[52]),
        .Q(R[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[60]),
        .Q(R[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[2]),
        .Q(R[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[10]),
        .Q(R[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[18]),
        .Q(R[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[6]),
        .Q(R[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[26]),
        .Q(R[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[34]),
        .Q(R[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[42]),
        .Q(R[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[50]),
        .Q(R[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[58]),
        .Q(R[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[0]),
        .Q(R[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[8]),
        .Q(R[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[16]),
        .Q(R[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[24]),
        .Q(R[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[32]),
        .Q(R[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[14]),
        .Q(R[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[40]),
        .Q(R[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[48]),
        .Q(R[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[56]),
        .Q(R[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[22]),
        .Q(R[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[30]),
        .Q(R[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[38]),
        .Q(R[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[46]),
        .Q(R[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[54]),
        .Q(R[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[62]),
        .Q(R[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \R_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desOut[4]),
        .Q(R[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC
       (.P(\<const1>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[0]_INST_0 
       (.I0(desIn[0]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[25]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[57] ),
        .I5(out[25]),
        .O(desOut[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[10]_INST_0 
       (.I0(desIn[10]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[18]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[50] ),
        .I5(out[18]),
        .O(desOut[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[11]_INST_0 
       (.I0(R[18]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[50] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[11]),
        .O(desOut[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[12]_INST_0 
       (.I0(desIn[12]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[10]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[42] ),
        .I5(out[10]),
        .O(desOut[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[13]_INST_0 
       (.I0(R[10]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[42] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[13]),
        .O(desOut[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[14]_INST_0 
       (.I0(desIn[14]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[2]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[34] ),
        .I5(out[2]),
        .O(desOut[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[15]_INST_0 
       (.I0(R[2]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[34] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[15]),
        .O(desOut[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[16]_INST_0 
       (.I0(desIn[16]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[27]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[59] ),
        .I5(out[27]),
        .O(desOut[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[17]_INST_0 
       (.I0(R[27]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[59] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[17]),
        .O(desOut[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[18]_INST_0 
       (.I0(desIn[18]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[19]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[51] ),
        .I5(out[19]),
        .O(desOut[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[19]_INST_0 
       (.I0(R[19]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[51] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[19]),
        .O(desOut[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[1]_INST_0 
       (.I0(R[25]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[57] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[1]),
        .O(desOut[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[20]_INST_0 
       (.I0(desIn[20]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[11]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[43] ),
        .I5(out[11]),
        .O(desOut[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[21]_INST_0 
       (.I0(R[11]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[43] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[21]),
        .O(desOut[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[22]_INST_0 
       (.I0(desIn[22]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[3]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[35] ),
        .I5(out[3]),
        .O(desOut[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[23]_INST_0 
       (.I0(R[3]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[35] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[23]),
        .O(desOut[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[24]_INST_0 
       (.I0(desIn[24]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[28]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[60] ),
        .I5(out[28]),
        .O(desOut[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[25]_INST_0 
       (.I0(R[28]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[60] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[25]),
        .O(desOut[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[26]_INST_0 
       (.I0(desIn[26]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[20]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[52] ),
        .I5(out[20]),
        .O(desOut[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[27]_INST_0 
       (.I0(R[20]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[52] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[27]),
        .O(desOut[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[28]_INST_0 
       (.I0(desIn[28]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[12]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[44] ),
        .I5(out[12]),
        .O(desOut[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[29]_INST_0 
       (.I0(R[12]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[44] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[29]),
        .O(desOut[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[2]_INST_0 
       (.I0(desIn[2]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[17]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[49] ),
        .I5(out[17]),
        .O(desOut[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[30]_INST_0 
       (.I0(desIn[30]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[4]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[36] ),
        .I5(out[4]),
        .O(desOut[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[31]_INST_0 
       (.I0(R[4]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[36] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[31]),
        .O(desOut[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[32]_INST_0 
       (.I0(desIn[32]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[29]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[61] ),
        .I5(out[29]),
        .O(desOut[32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[33]_INST_0 
       (.I0(R[29]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[61] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[33]),
        .O(desOut[33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[34]_INST_0 
       (.I0(desIn[34]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[21]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[53] ),
        .I5(out[21]),
        .O(desOut[34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[35]_INST_0 
       (.I0(R[21]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[53] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[35]),
        .O(desOut[35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[36]_INST_0 
       (.I0(desIn[36]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[13]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[45] ),
        .I5(out[13]),
        .O(desOut[36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[37]_INST_0 
       (.I0(R[13]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[45] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[37]),
        .O(desOut[37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[38]_INST_0 
       (.I0(desIn[38]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[5]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[37] ),
        .I5(out[5]),
        .O(desOut[38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[39]_INST_0 
       (.I0(R[5]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[37] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[39]),
        .O(desOut[39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[3]_INST_0 
       (.I0(R[17]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[49] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[3]),
        .O(desOut[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[40]_INST_0 
       (.I0(desIn[40]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[30]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[62] ),
        .I5(out[30]),
        .O(desOut[40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[41]_INST_0 
       (.I0(R[30]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[62] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[41]),
        .O(desOut[41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[42]_INST_0 
       (.I0(desIn[42]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[22]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[54] ),
        .I5(out[22]),
        .O(desOut[42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[43]_INST_0 
       (.I0(R[22]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[54] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[43]),
        .O(desOut[43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[44]_INST_0 
       (.I0(desIn[44]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[14]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[46] ),
        .I5(out[14]),
        .O(desOut[44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[45]_INST_0 
       (.I0(R[14]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[46] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[45]),
        .O(desOut[45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[46]_INST_0 
       (.I0(desIn[46]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[6]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[38] ),
        .I5(out[6]),
        .O(desOut[46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[47]_INST_0 
       (.I0(R[6]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[38] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[47]),
        .O(desOut[47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[48]_INST_0 
       (.I0(desIn[48]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[31]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[63] ),
        .I5(out[31]),
        .O(desOut[48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[49]_INST_0 
       (.I0(R[31]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[63] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[49]),
        .O(desOut[49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[4]_INST_0 
       (.I0(desIn[4]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[9]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[41] ),
        .I5(out[9]),
        .O(desOut[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[50]_INST_0 
       (.I0(desIn[50]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[23]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[55] ),
        .I5(out[23]),
        .O(desOut[50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[51]_INST_0 
       (.I0(R[23]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[55] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[51]),
        .O(desOut[51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[52]_INST_0 
       (.I0(desIn[52]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[15]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[47] ),
        .I5(out[15]),
        .O(desOut[52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[53]_INST_0 
       (.I0(R[15]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[47] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[53]),
        .O(desOut[53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[54]_INST_0 
       (.I0(desIn[54]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[7]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[39] ),
        .I5(out[7]),
        .O(desOut[54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[55]_INST_0 
       (.I0(R[7]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[39] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[55]),
        .O(desOut[55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[56]_INST_0 
       (.I0(desIn[56]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[32]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[64] ),
        .I5(out[32]),
        .O(desOut[56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[57]_INST_0 
       (.I0(R[32]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[64] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[57]),
        .O(desOut[57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[58]_INST_0 
       (.I0(desIn[58]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[24]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[56] ),
        .I5(out[24]),
        .O(desOut[58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[59]_INST_0 
       (.I0(R[24]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[56] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[59]),
        .O(desOut[59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[5]_INST_0 
       (.I0(R[9]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[41] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[5]),
        .O(desOut[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[60]_INST_0 
       (.I0(desIn[60]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[16]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[48] ),
        .I5(out[16]),
        .O(desOut[60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[61]_INST_0 
       (.I0(R[16]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[48] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[61]),
        .O(desOut[61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[62]_INST_0 
       (.I0(desIn[62]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[8]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[40] ),
        .I5(out[8]),
        .O(desOut[62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \desOut[62]_INST_0_i_1 
       (.I0(roundSel[4]),
        .I1(roundSel[5]),
        .O(\desOut[62]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \desOut[62]_INST_0_i_2 
       (.I0(roundSel[0]),
        .I1(roundSel[1]),
        .I2(roundSel[5]),
        .I3(roundSel[4]),
        .I4(roundSel[3]),
        .I5(roundSel[2]),
        .O(\desOut[62]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[63]_INST_0 
       (.I0(R[8]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[40] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[63]),
        .O(desOut[63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEF)) 
    \desOut[63]_INST_0_i_1 
       (.I0(roundSel[3]),
        .I1(roundSel[1]),
        .I2(roundSel[5]),
        .I3(roundSel[4]),
        .I4(roundSel[0]),
        .I5(roundSel[2]),
        .O(\desOut[63]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \desOut[63]_INST_0_i_2 
       (.I0(roundSel[5]),
        .I1(roundSel[4]),
        .I2(roundSel[1]),
        .I3(roundSel[0]),
        .I4(roundSel[3]),
        .I5(roundSel[2]),
        .O(\desOut[63]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[6]_INST_0 
       (.I0(desIn[6]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[1]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(FP_R_reg_n_0_),
        .I5(out[1]),
        .O(desOut[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[7]_INST_0 
       (.I0(R[1]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(FP_R_reg_n_0_),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[7]),
        .O(desOut[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001DFF1DFFE200E2)) 
    \desOut[8]_INST_0 
       (.I0(desIn[8]),
        .I1(\desOut[62]_INST_0_i_1_n_0 ),
        .I2(R[26]),
        .I3(\desOut[62]_INST_0_i_2_n_0 ),
        .I4(\FP_R_reg_n_0_[58] ),
        .I5(out[26]),
        .O(desOut[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \desOut[9]_INST_0 
       (.I0(R[26]),
        .I1(\desOut[63]_INST_0_i_1_n_0 ),
        .I2(\FP_R_reg_n_0_[58] ),
        .I3(\desOut[63]_INST_0_i_2_n_0 ),
        .I4(desIn[9]),
        .O(desOut[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0
       (.I0(\u0/X [41]),
        .I1(\u0/X [40]),
        .I2(\u0/X [39]),
        .I3(\u0/X [38]),
        .I4(\u0/X [42]),
        .I5(\u0/X [37]),
        .O(out[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__0
       (.I0(\u0/X [17]),
        .I1(\u0/X [16]),
        .I2(\u0/X [15]),
        .I3(\u0/X [14]),
        .I4(\u0/X [18]),
        .I5(\u0/X [13]),
        .O(out[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__1
       (.I0(\u0/X [35]),
        .I1(\u0/X [34]),
        .I2(\u0/X [33]),
        .I3(\u0/X [32]),
        .I4(\u0/X [36]),
        .I5(\u0/X [31]),
        .O(out[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__2
       (.I0(\u0/X [11]),
        .I1(\u0/X [10]),
        .I2(\u0/X [9]),
        .I3(\u0/X [8]),
        .I4(\u0/X [12]),
        .I5(\u0/X [7]),
        .O(out[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__3
       (.I0(\u0/X [47]),
        .I1(\u0/X [46]),
        .I2(\u0/X [45]),
        .I3(\u0/X [44]),
        .I4(\u0/X [48]),
        .I5(\u0/X [43]),
        .O(out[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__4
       (.I0(\u0/X [23]),
        .I1(\u0/X [22]),
        .I2(\u0/X [21]),
        .I3(\u0/X [20]),
        .I4(\u0/X [24]),
        .I5(\u0/X [19]),
        .O(out[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__5
       (.I0(\u0/X [29]),
        .I1(\u0/X [28]),
        .I2(\u0/X [27]),
        .I3(\u0/X [26]),
        .I4(\u0/X [30]),
        .I5(\u0/X [25]),
        .O(out[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__6
       (.I0(\u0/X [5]),
        .I1(\u0/X [4]),
        .I2(\u0/X [3]),
        .I3(\u0/X [2]),
        .I4(\u0/X [6]),
        .I5(\u0/X [1]),
        .O(out[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_1
       (.I0(desOut[25]),
        .I1(g0_b0_i_7_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_8_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_9_n_0),
        .O(\u0/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_10
       (.I0(g0_b0_i_31_n_0),
        .I1(g0_b0_i_32__6_n_0),
        .O(g0_b0_i_10_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_100
       (.I0(g0_b0_i_124_n_0),
        .I1(\u1/decrypt_int__2 ),
        .I2(g0_b0_i_99__1_n_0),
        .O(g0_b0_i_100_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_100__0
       (.I0(key3[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_65__4_n_0),
        .I3(roundSel[4]),
        .I4(key1[0]),
        .O(g0_b0_i_100__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_100__1
       (.I0(key2[7]),
        .I1(roundSel[5]),
        .I2(key3[7]),
        .I3(decrypt),
        .I4(key1[7]),
        .I5(roundSel[4]),
        .O(g0_b0_i_100__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_100__2
       (.I0(key2[19]),
        .I1(roundSel[5]),
        .I2(key3[19]),
        .I3(decrypt),
        .I4(key1[19]),
        .I5(roundSel[4]),
        .O(\u1/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_101
       (.I0(\u1/p_2_in ),
        .I1(\u1/p_3_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_16_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_96__2_n_0),
        .O(g0_b0_i_101_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_101__0
       (.I0(g0_b0_i_67__5_n_0),
        .I1(\u1/decrypt_int__2 ),
        .I2(g0_b0_i_71__5_n_0),
        .O(g0_b0_i_101__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_101__1
       (.I0(g0_b0_i_71__5_n_0),
        .I1(\u1/decrypt_int__2 ),
        .I2(g0_b0_i_88__3_n_0),
        .O(g0_b0_i_101__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_101__2
       (.I0(key2[15]),
        .I1(roundSel[5]),
        .I2(key3[15]),
        .I3(decrypt),
        .I4(key1[15]),
        .I5(roundSel[4]),
        .O(g0_b0_i_101__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_102
       (.I0(\u1/p_1_in ),
        .I1(\u1/p_14_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_19_in ),
        .I4(g0_b0_i_74__6_n_0),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_102_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_102__0
       (.I0(g0_b0_i_71__5_n_0),
        .I1(\u1/decrypt_int__2 ),
        .I2(g0_b0_i_99__1_n_0),
        .O(g0_b0_i_102__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_102__1
       (.I0(key1[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_79__6_n_0),
        .I3(roundSel[4]),
        .I4(key3[0]),
        .O(g0_b0_i_102__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_102__2
       (.I0(key2[29]),
        .I1(roundSel[5]),
        .I2(key3[29]),
        .I3(decrypt),
        .I4(key1[29]),
        .I5(roundSel[4]),
        .O(g0_b0_i_102__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_103
       (.I0(g0_b0_i_67__5_n_0),
        .I1(g0_b0_i_66__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_69__5_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_110__0_n_0),
        .O(g0_b0_i_103_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_103__0
       (.I0(\u1/p_17_in ),
        .I1(\u1/p_9_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_67__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_77__5_n_0),
        .O(g0_b0_i_103__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_103__1
       (.I0(key1[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_119_n_0),
        .I3(roundSel[4]),
        .I4(key3[0]),
        .O(g0_b0_i_103__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_104
       (.I0(g0_b0_i_72__6_n_0),
        .I1(g0_b0_i_71__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_65__4_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_73__6_n_0),
        .O(g0_b0_i_104_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_104__0
       (.I0(\u1/p_7_in ),
        .I1(g0_b0_i_89__3_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_71__6_n_0),
        .I4(\u1/p_10_in ),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_104__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_104__1
       (.I0(key1[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_90__3_n_0),
        .I3(roundSel[4]),
        .I4(key3[0]),
        .O(g0_b0_i_104__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_105
       (.I0(g0_b0_i_100__1_n_0),
        .I1(\u1/decrypt_int__2 ),
        .I2(g0_b0_i_124_n_0),
        .O(g0_b0_i_105_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_105__0
       (.I0(\u1/p_13_in ),
        .I1(\u1/p_17_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_71__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_98__1_n_0),
        .O(g0_b0_i_105__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_105__1
       (.I0(g0_b0_i_128_n_0),
        .I1(roundSel[0]),
        .I2(g0_b0_i_108__0_n_0),
        .I3(decrypt),
        .I4(g0_b0_i_129_n_0),
        .O(g0_b0_i_105__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_106
       (.I0(\u1/p_10_in ),
        .I1(\u1/p_1_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_89__3_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_67__6_n_0),
        .O(g0_b0_i_106_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_106__0
       (.I0(g0_b0_i_79__6_n_0),
        .I1(g0_b0_i_77__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_88__3_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_80__6_n_0),
        .O(g0_b0_i_106__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_107
       (.I0(g0_b0_i_77__5_n_0),
        .I1(\u1/p_2_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_9_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_19_in ),
        .O(g0_b0_i_107_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_107__0
       (.I0(key1[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_70__6_n_0),
        .I3(roundSel[4]),
        .I4(key3[0]),
        .O(g0_b0_i_107__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_108
       (.I0(g0_b0_i_74__6_n_0),
        .I1(\u1/p_15_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_14_in ),
        .I4(g0_b0_i_96__2_n_0),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_108_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFB08)) 
    g0_b0_i_108__0
       (.I0(key2[0]),
        .I1(roundSel[4]),
        .I2(roundSel[5]),
        .I3(g0_b0_i_70__6_n_0),
        .O(g0_b0_i_108__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_109
       (.I0(\u1/p_15_in ),
        .I1(\u1/p_14_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_74__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_95__2_n_0),
        .O(g0_b0_i_109_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_109__0
       (.I0(g0_b0_i_124_n_0),
        .I1(g0_b0_i_68__6_n_0),
        .I2(g0_b0_i_85__3_n_0),
        .O(g0_b0_i_109__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_10__0
       (.I0(g0_b0_i_31__0_n_0),
        .I1(g0_b0_i_32__0_n_0),
        .O(g0_b0_i_10__0_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_10__1
       (.I0(g0_b0_i_31__1_n_0),
        .I1(g0_b0_i_32__1_n_0),
        .O(g0_b0_i_10__1_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_10__2
       (.I0(g0_b0_i_31__2_n_0),
        .I1(g0_b0_i_32__2_n_0),
        .O(g0_b0_i_10__2_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_10__3
       (.I0(g0_b0_i_31__3_n_0),
        .I1(g0_b0_i_32__3_n_0),
        .O(g0_b0_i_10__3_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_10__4
       (.I0(g0_b0_i_31__4_n_0),
        .I1(g0_b0_i_32__4_n_0),
        .O(g0_b0_i_10__4_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_10__5
       (.I0(g0_b0_i_31__5_n_0),
        .I1(g0_b0_i_32__5_n_0),
        .O(g0_b0_i_10__5_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_10__6
       (.I0(g0_b0_i_31__6_n_0),
        .I1(g0_b0_i_32_n_0),
        .O(g0_b0_i_10__6_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_11
       (.I0(g0_b0_i_33_n_0),
        .I1(g0_b0_i_34_n_0),
        .O(g0_b0_i_11_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_110
       (.I0(\u1/p_2_in ),
        .I1(\u1/p_9_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_96__2_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_77__5_n_0),
        .O(g0_b0_i_110_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_110__0
       (.I0(key2[37]),
        .I1(roundSel[5]),
        .I2(key3[37]),
        .I3(decrypt),
        .I4(key1[37]),
        .I5(roundSel[4]),
        .O(g0_b0_i_110__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_111
       (.I0(g0_b0_i_119_n_0),
        .I1(g0_b0_i_71__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_73__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_99__1_n_0),
        .O(g0_b0_i_111_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_111__0
       (.I0(\u1/p_1_in ),
        .I1(g0_b0_i_89__3_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_19_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_10_in ),
        .O(g0_b0_i_111__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_112
       (.I0(g0_b0_i_130_n_0),
        .I1(roundSel[0]),
        .I2(g0_b0_i_117_n_0),
        .I3(decrypt),
        .I4(g0_b0_i_131_n_0),
        .O(g0_b0_i_112_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_112__0
       (.I0(\u1/p_17_in ),
        .I1(g0_b0_i_98__1_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_67__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_13_in ),
        .O(g0_b0_i_112__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_113
       (.I0(g0_b0_i_72__6_n_0),
        .I1(g0_b0_i_77__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_65__4_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_80__6_n_0),
        .O(g0_b0_i_113_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_114
       (.I0(g0_b0_i_85__3_n_0),
        .I1(g0_b0_i_101__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_70__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_115_n_0),
        .O(g0_b0_i_114_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_115
       (.I0(key2[1]),
        .I1(roundSel[5]),
        .I2(key3[1]),
        .I3(decrypt),
        .I4(key1[1]),
        .I5(roundSel[4]),
        .O(g0_b0_i_115_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_116
       (.I0(key1[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_110__0_n_0),
        .I3(roundSel[4]),
        .I4(key3[0]),
        .O(g0_b0_i_116_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFB08)) 
    g0_b0_i_117
       (.I0(key2[0]),
        .I1(roundSel[4]),
        .I2(roundSel[5]),
        .I3(g0_b0_i_110__0_n_0),
        .O(g0_b0_i_117_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_118
       (.I0(g0_b0_i_124_n_0),
        .I1(g0_b0_i_68__6_n_0),
        .I2(g0_b0_i_67__5_n_0),
        .O(g0_b0_i_118_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_119
       (.I0(key2[51]),
        .I1(roundSel[5]),
        .I2(key3[51]),
        .I3(decrypt),
        .I4(key1[51]),
        .I5(roundSel[4]),
        .O(g0_b0_i_119_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_11__0
       (.I0(g0_b0_i_33__0_n_0),
        .I1(g0_b0_i_34__0_n_0),
        .O(g0_b0_i_11__0_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_11__1
       (.I0(g0_b0_i_33__1_n_0),
        .I1(g0_b0_i_34__2_n_0),
        .O(g0_b0_i_11__1_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_11__2
       (.I0(g0_b0_i_33__2_n_0),
        .I1(g0_b0_i_34__1_n_0),
        .O(g0_b0_i_11__2_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_11__3
       (.I0(g0_b0_i_33__3_n_0),
        .I1(g0_b0_i_34__5_n_0),
        .O(g0_b0_i_11__3_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_11__4
       (.I0(g0_b0_i_33__4_n_0),
        .I1(g0_b0_i_34__6_n_0),
        .O(g0_b0_i_11__4_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_11__5
       (.I0(g0_b0_i_33__5_n_0),
        .I1(g0_b0_i_34__3_n_0),
        .O(g0_b0_i_11__5_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_11__6
       (.I0(g0_b0_i_33__6_n_0),
        .I1(g0_b0_i_34__4_n_0),
        .O(g0_b0_i_11__6_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_12
       (.I0(g0_b0_i_35_n_0),
        .I1(g0_b0_i_36_n_0),
        .O(g0_b0_i_12_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_120
       (.I0(g0_b0_i_87__3_n_0),
        .I1(g0_b0_i_65__4_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_72__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_86__2_n_0),
        .O(g0_b0_i_120_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_121
       (.I0(g0_b0_i_101__2_n_0),
        .I1(g0_b0_i_110__0_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_102__2_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_67__5_n_0),
        .O(g0_b0_i_121_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_122
       (.I0(g0_b0_i_77__6_n_0),
        .I1(g0_b0_i_99__1_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_115_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_119_n_0),
        .O(g0_b0_i_122_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_123
       (.I0(g0_b0_i_124_n_0),
        .I1(g0_b0_i_100__1_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_80__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_98__2_n_0),
        .O(g0_b0_i_123_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_124
       (.I0(key2[14]),
        .I1(roundSel[5]),
        .I2(key3[14]),
        .I3(decrypt),
        .I4(key1[14]),
        .I5(roundSel[4]),
        .O(g0_b0_i_124_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_125
       (.I0(key1[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_85__3_n_0),
        .I3(roundSel[4]),
        .I4(key3[0]),
        .O(g0_b0_i_125_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_126
       (.I0(g0_b0_i_124_n_0),
        .I1(g0_b0_i_68__6_n_0),
        .I2(g0_b0_i_88__3_n_0),
        .O(g0_b0_i_126_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_127
       (.I0(g0_b0_i_71__5_n_0),
        .I1(g0_b0_i_68__6_n_0),
        .I2(g0_b0_i_100__1_n_0),
        .O(g0_b0_i_127_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_128
       (.I0(g0_b0_i_85__3_n_0),
        .I1(g0_b0_i_68__6_n_0),
        .I2(g0_b0_i_124_n_0),
        .O(g0_b0_i_128_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_129
       (.I0(key3[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_70__6_n_0),
        .I3(roundSel[4]),
        .I4(key1[0]),
        .O(g0_b0_i_129_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_12__0
       (.I0(g0_b0_i_35__2_n_0),
        .I1(g0_b0_i_36__0_n_0),
        .O(g0_b0_i_12__0_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_12__1
       (.I0(g0_b0_i_35__1_n_0),
        .I1(g0_b0_i_36__1_n_0),
        .O(g0_b0_i_12__1_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_12__2
       (.I0(g0_b0_i_35__4_n_0),
        .I1(g0_b0_i_36__2_n_0),
        .O(g0_b0_i_12__2_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_12__3
       (.I0(g0_b0_i_35__5_n_0),
        .I1(g0_b0_i_36__3_n_0),
        .O(g0_b0_i_12__3_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_12__4
       (.I0(g0_b0_i_35__6_n_0),
        .I1(g0_b0_i_36__4_n_0),
        .O(g0_b0_i_12__4_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_12__5
       (.I0(g0_b0_i_35__0_n_0),
        .I1(g0_b0_i_36__5_n_0),
        .O(g0_b0_i_12__5_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_12__6
       (.I0(g0_b0_i_35__3_n_0),
        .I1(g0_b0_i_36__6_n_0),
        .O(g0_b0_i_12__6_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_13
       (.I0(g0_b0_i_37_n_0),
        .I1(g0_b0_i_38_n_0),
        .O(g0_b0_i_13_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_130
       (.I0(g0_b0_i_67__5_n_0),
        .I1(g0_b0_i_68__6_n_0),
        .I2(g0_b0_i_124_n_0),
        .O(g0_b0_i_130_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_131
       (.I0(key3[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_110__0_n_0),
        .I3(roundSel[4]),
        .I4(key1[0]),
        .O(g0_b0_i_131_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_13__0
       (.I0(g0_b0_i_37__0_n_0),
        .I1(g0_b0_i_38__0_n_0),
        .O(g0_b0_i_13__0_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_13__1
       (.I0(g0_b0_i_37__1_n_0),
        .I1(g0_b0_i_38__1_n_0),
        .O(g0_b0_i_13__1_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_13__2
       (.I0(g0_b0_i_37__2_n_0),
        .I1(g0_b0_i_38__2_n_0),
        .O(g0_b0_i_13__2_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_13__3
       (.I0(g0_b0_i_37__3_n_0),
        .I1(g0_b0_i_38__5_n_0),
        .O(g0_b0_i_13__3_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_13__4
       (.I0(g0_b0_i_37__4_n_0),
        .I1(g0_b0_i_38__6_n_0),
        .O(g0_b0_i_13__4_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_13__5
       (.I0(g0_b0_i_37__5_n_0),
        .I1(g0_b0_i_38__3_n_0),
        .O(g0_b0_i_13__5_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_13__6
       (.I0(g0_b0_i_37__6_n_0),
        .I1(g0_b0_i_38__4_n_0),
        .O(g0_b0_i_13__6_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_14
       (.I0(g0_b0_i_39_n_0),
        .I1(g0_b0_i_40_n_0),
        .O(g0_b0_i_14_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_14__0
       (.I0(g0_b0_i_39__0_n_0),
        .I1(g0_b0_i_40__0_n_0),
        .O(g0_b0_i_14__0_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_14__1
       (.I0(g0_b0_i_39__1_n_0),
        .I1(g0_b0_i_40__2_n_0),
        .O(g0_b0_i_14__1_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_14__2
       (.I0(g0_b0_i_39__2_n_0),
        .I1(g0_b0_i_40__1_n_0),
        .O(g0_b0_i_14__2_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_14__3
       (.I0(g0_b0_i_39__3_n_0),
        .I1(g0_b0_i_40__3_n_0),
        .O(g0_b0_i_14__3_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_14__4
       (.I0(g0_b0_i_39__4_n_0),
        .I1(g0_b0_i_40__4_n_0),
        .O(g0_b0_i_14__4_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_14__5
       (.I0(g0_b0_i_39__5_n_0),
        .I1(g0_b0_i_40__6_n_0),
        .O(g0_b0_i_14__5_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_14__6
       (.I0(g0_b0_i_39__6_n_0),
        .I1(g0_b0_i_40__5_n_0),
        .O(g0_b0_i_14__6_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_15
       (.I0(g0_b0_i_41_n_0),
        .I1(g0_b0_i_42_n_0),
        .O(g0_b0_i_15_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_15__0
       (.I0(g0_b0_i_41__0_n_0),
        .I1(g0_b0_i_42__0_n_0),
        .O(g0_b0_i_15__0_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_15__1
       (.I0(g0_b0_i_41__1_n_0),
        .I1(g0_b0_i_42__1_n_0),
        .O(g0_b0_i_15__1_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_15__2
       (.I0(g0_b0_i_41__6_n_0),
        .I1(g0_b0_i_42__2_n_0),
        .O(g0_b0_i_15__2_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_15__3
       (.I0(g0_b0_i_41__2_n_0),
        .I1(g0_b0_i_42__3_n_0),
        .O(g0_b0_i_15__3_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_15__4
       (.I0(g0_b0_i_41__3_n_0),
        .I1(g0_b0_i_42__4_n_0),
        .O(g0_b0_i_15__4_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_15__5
       (.I0(g0_b0_i_41__4_n_0),
        .I1(g0_b0_i_42__5_n_0),
        .O(g0_b0_i_15__5_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_15__6
       (.I0(g0_b0_i_41__5_n_0),
        .I1(g0_b0_i_42__6_n_0),
        .O(g0_b0_i_15__6_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_16
       (.I0(g0_b0_i_43_n_0),
        .I1(g0_b0_i_44_n_0),
        .O(g0_b0_i_16_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_16__0
       (.I0(g0_b0_i_43__0_n_0),
        .I1(g0_b0_i_44__6_n_0),
        .O(g0_b0_i_16__0_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_16__1
       (.I0(g0_b0_i_43__1_n_0),
        .I1(g0_b0_i_44__0_n_0),
        .O(g0_b0_i_16__1_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_16__2
       (.I0(g0_b0_i_43__2_n_0),
        .I1(g0_b0_i_44__1_n_0),
        .O(g0_b0_i_16__2_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_16__3
       (.I0(g0_b0_i_43__3_n_0),
        .I1(g0_b0_i_44__2_n_0),
        .O(g0_b0_i_16__3_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_16__4
       (.I0(g0_b0_i_43__4_n_0),
        .I1(g0_b0_i_44__3_n_0),
        .O(g0_b0_i_16__4_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_16__5
       (.I0(g0_b0_i_43__5_n_0),
        .I1(g0_b0_i_44__4_n_0),
        .O(g0_b0_i_16__5_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_16__6
       (.I0(g0_b0_i_43__6_n_0),
        .I1(g0_b0_i_44__5_n_0),
        .O(g0_b0_i_16__6_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_17
       (.I0(g0_b0_i_45_n_0),
        .I1(g0_b0_i_46__3_n_0),
        .O(g0_b0_i_17_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_17__0
       (.I0(g0_b0_i_45__0_n_0),
        .I1(g0_b0_i_46__6_n_0),
        .O(g0_b0_i_17__0_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_17__1
       (.I0(g0_b0_i_45__1_n_0),
        .I1(g0_b0_i_46__4_n_0),
        .O(g0_b0_i_17__1_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_17__2
       (.I0(g0_b0_i_45__2_n_0),
        .I1(g0_b0_i_46__5_n_0),
        .O(g0_b0_i_17__2_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_17__3
       (.I0(g0_b0_i_45__3_n_0),
        .I1(g0_b0_i_46__0_n_0),
        .O(g0_b0_i_17__3_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_17__4
       (.I0(g0_b0_i_45__4_n_0),
        .I1(g0_b0_i_46__1_n_0),
        .O(g0_b0_i_17__4_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_17__5
       (.I0(g0_b0_i_45__5_n_0),
        .I1(g0_b0_i_46__2_n_0),
        .O(g0_b0_i_17__5_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_17__6
       (.I0(g0_b0_i_45__6_n_0),
        .I1(g0_b0_i_46_n_0),
        .O(g0_b0_i_17__6_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_18
       (.I0(g0_b0_i_47_n_0),
        .I1(g0_b0_i_48_n_0),
        .O(g0_b0_i_18_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_18__0
       (.I0(g0_b0_i_47__3_n_0),
        .I1(g0_b0_i_48__0_n_0),
        .O(g0_b0_i_18__0_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_18__1
       (.I0(g0_b0_i_47__6_n_0),
        .I1(g0_b0_i_48__1_n_0),
        .O(g0_b0_i_18__1_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_18__2
       (.I0(g0_b0_i_47__4_n_0),
        .I1(g0_b0_i_48__2_n_0),
        .O(g0_b0_i_18__2_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_18__3
       (.I0(g0_b0_i_47__5_n_0),
        .I1(g0_b0_i_48__3_n_0),
        .O(g0_b0_i_18__3_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_18__4
       (.I0(g0_b0_i_47__0_n_0),
        .I1(g0_b0_i_48__4_n_0),
        .O(g0_b0_i_18__4_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_18__5
       (.I0(g0_b0_i_47__1_n_0),
        .I1(g0_b0_i_48__5_n_0),
        .O(g0_b0_i_18__5_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_18__6
       (.I0(g0_b0_i_47__2_n_0),
        .I1(g0_b0_i_48__6_n_0),
        .O(g0_b0_i_18__6_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_19
       (.I0(g0_b0_i_49_n_0),
        .I1(g0_b0_i_50_n_0),
        .O(g0_b0_i_19_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_19__0
       (.I0(g0_b0_i_49__0_n_0),
        .I1(g0_b0_i_50__0_n_0),
        .O(g0_b0_i_19__0_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_19__1
       (.I0(g0_b0_i_49__1_n_0),
        .I1(g0_b0_i_50__1_n_0),
        .O(g0_b0_i_19__1_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_19__2
       (.I0(g0_b0_i_49__2_n_0),
        .I1(g0_b0_i_50__2_n_0),
        .O(g0_b0_i_19__2_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_19__3
       (.I0(g0_b0_i_49__3_n_0),
        .I1(g0_b0_i_50__3_n_0),
        .O(g0_b0_i_19__3_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_19__4
       (.I0(g0_b0_i_49__4_n_0),
        .I1(g0_b0_i_50__4_n_0),
        .O(g0_b0_i_19__4_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_19__5
       (.I0(g0_b0_i_49__5_n_0),
        .I1(g0_b0_i_50__5_n_0),
        .O(g0_b0_i_19__5_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_19__6
       (.I0(g0_b0_i_49__6_n_0),
        .I1(g0_b0_i_50__6_n_0),
        .O(g0_b0_i_19__6_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_1__0
       (.I0(desOut[59]),
        .I1(g0_b0_i_7__0_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_8__1_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_9__1_n_0),
        .O(\u0/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_1__1
       (.I0(desOut[27]),
        .I1(g0_b0_i_7__1_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_8__0_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_9__0_n_0),
        .O(\u0/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_1__2
       (.I0(desOut[61]),
        .I1(g0_b0_i_7__2_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_8__2_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_9__2_n_0),
        .O(\u0/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_1__3
       (.I0(desOut[63]),
        .I1(g0_b0_i_7__4_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_8__3_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_9__3_n_0),
        .O(\u0/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_1__4
       (.I0(desOut[29]),
        .I1(g0_b0_i_7__3_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_8__4_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_9__4_n_0),
        .O(\u0/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_1__5
       (.I0(desOut[31]),
        .I1(g0_b0_i_7__5_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_8__5_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_9__5_n_0),
        .O(\u0/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_1__6
       (.I0(desOut[57]),
        .I1(g0_b0_i_7__6_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_8__6_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_9__6_n_0),
        .O(\u0/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_2
       (.I0(desOut[49]),
        .I1(g0_b0_i_10_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_11_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_12_n_0),
        .O(\u0/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_20
       (.I0(g0_b0_i_51_n_0),
        .I1(g0_b0_i_52_n_0),
        .O(g0_b0_i_20_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_20__0
       (.I0(g0_b0_i_51__0_n_0),
        .I1(g0_b0_i_52__1_n_0),
        .O(g0_b0_i_20__0_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_20__1
       (.I0(g0_b0_i_51__1_n_0),
        .I1(g0_b0_i_52__0_n_0),
        .O(g0_b0_i_20__1_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_20__2
       (.I0(g0_b0_i_51__2_n_0),
        .I1(g0_b0_i_52__2_n_0),
        .O(g0_b0_i_20__2_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_20__3
       (.I0(g0_b0_i_51__3_n_0),
        .I1(g0_b0_i_52__3_n_0),
        .O(g0_b0_i_20__3_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_20__4
       (.I0(g0_b0_i_51__4_n_0),
        .I1(g0_b0_i_52__6_n_0),
        .O(g0_b0_i_20__4_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_20__5
       (.I0(g0_b0_i_51__5_n_0),
        .I1(g0_b0_i_52__5_n_0),
        .O(g0_b0_i_20__5_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_20__6
       (.I0(g0_b0_i_51__6_n_0),
        .I1(g0_b0_i_52__4_n_0),
        .O(g0_b0_i_20__6_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_21
       (.I0(g0_b0_i_53_n_0),
        .I1(g0_b0_i_54_n_0),
        .O(g0_b0_i_21_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_21__0
       (.I0(g0_b0_i_53__1_n_0),
        .I1(g0_b0_i_54__0_n_0),
        .O(g0_b0_i_21__0_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_21__1
       (.I0(g0_b0_i_53__0_n_0),
        .I1(g0_b0_i_54__1_n_0),
        .O(g0_b0_i_21__1_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_21__2
       (.I0(g0_b0_i_53__2_n_0),
        .I1(g0_b0_i_54__2_n_0),
        .O(g0_b0_i_21__2_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_21__3
       (.I0(g0_b0_i_53__3_n_0),
        .I1(g0_b0_i_54__3_n_0),
        .O(g0_b0_i_21__3_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_21__4
       (.I0(g0_b0_i_53__6_n_0),
        .I1(g0_b0_i_54__4_n_0),
        .O(g0_b0_i_21__4_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_21__5
       (.I0(g0_b0_i_53__5_n_0),
        .I1(g0_b0_i_54__5_n_0),
        .O(g0_b0_i_21__5_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_21__6
       (.I0(g0_b0_i_53__4_n_0),
        .I1(g0_b0_i_54__6_n_0),
        .O(g0_b0_i_21__6_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_22
       (.I0(g0_b0_i_55_n_0),
        .I1(g0_b0_i_56_n_0),
        .O(g0_b0_i_22_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_22__0
       (.I0(g0_b0_i_55__0_n_0),
        .I1(g0_b0_i_56__0_n_0),
        .O(g0_b0_i_22__0_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_22__1
       (.I0(g0_b0_i_55__1_n_0),
        .I1(g0_b0_i_56__1_n_0),
        .O(g0_b0_i_22__1_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_22__2
       (.I0(g0_b0_i_55__2_n_0),
        .I1(g0_b0_i_56__2_n_0),
        .O(g0_b0_i_22__2_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_22__3
       (.I0(g0_b0_i_55__3_n_0),
        .I1(g0_b0_i_56__4_n_0),
        .O(g0_b0_i_22__3_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_22__4
       (.I0(g0_b0_i_55__4_n_0),
        .I1(g0_b0_i_56__3_n_0),
        .O(g0_b0_i_22__4_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_22__5
       (.I0(g0_b0_i_55__5_n_0),
        .I1(g0_b0_i_56__5_n_0),
        .O(g0_b0_i_22__5_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_22__6
       (.I0(g0_b0_i_55__6_n_0),
        .I1(g0_b0_i_56__6_n_0),
        .O(g0_b0_i_22__6_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_23
       (.I0(g0_b0_i_57_n_0),
        .I1(g0_b0_i_58_n_0),
        .O(g0_b0_i_23_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_23__0
       (.I0(g0_b0_i_57__0_n_0),
        .I1(g0_b0_i_58__1_n_0),
        .O(g0_b0_i_23__0_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_23__1
       (.I0(g0_b0_i_57__1_n_0),
        .I1(g0_b0_i_58__0_n_0),
        .O(g0_b0_i_23__1_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_23__2
       (.I0(g0_b0_i_57__2_n_0),
        .I1(g0_b0_i_58__2_n_0),
        .O(g0_b0_i_23__2_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_23__3
       (.I0(g0_b0_i_57__3_n_0),
        .I1(g0_b0_i_58__3_n_0),
        .O(g0_b0_i_23__3_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_23__4
       (.I0(g0_b0_i_57__4_n_0),
        .I1(g0_b0_i_58__6_n_0),
        .O(g0_b0_i_23__4_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_23__5
       (.I0(g0_b0_i_57__5_n_0),
        .I1(g0_b0_i_58__4_n_0),
        .O(g0_b0_i_23__5_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_23__6
       (.I0(g0_b0_i_57__6_n_0),
        .I1(g0_b0_i_58__5_n_0),
        .O(g0_b0_i_23__6_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_24
       (.I0(g0_b0_i_59_n_0),
        .I1(g0_b0_i_60_n_0),
        .O(g0_b0_i_24_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_24__0
       (.I0(g0_b0_i_59__1_n_0),
        .I1(g0_b0_i_60__0_n_0),
        .O(g0_b0_i_24__0_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_24__1
       (.I0(g0_b0_i_59__0_n_0),
        .I1(g0_b0_i_60__1_n_0),
        .O(g0_b0_i_24__1_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_24__2
       (.I0(g0_b0_i_59__2_n_0),
        .I1(g0_b0_i_60__2_n_0),
        .O(g0_b0_i_24__2_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_24__3
       (.I0(g0_b0_i_59__3_n_0),
        .I1(g0_b0_i_60__3_n_0),
        .O(g0_b0_i_24__3_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_24__4
       (.I0(g0_b0_i_59__6_n_0),
        .I1(g0_b0_i_60__4_n_0),
        .O(g0_b0_i_24__4_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_24__5
       (.I0(g0_b0_i_59__5_n_0),
        .I1(g0_b0_i_60__5_n_0),
        .O(g0_b0_i_24__5_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_24__6
       (.I0(g0_b0_i_59__4_n_0),
        .I1(g0_b0_i_60__6_n_0),
        .O(g0_b0_i_24__6_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_25
       (.I0(g0_b0_i_61_n_0),
        .I1(g0_b0_i_62__0_n_0),
        .O(g0_b0_i_25_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_25__0
       (.I0(g0_b0_i_61__0_n_0),
        .I1(g0_b0_i_62__1_n_0),
        .O(g0_b0_i_25__0_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_25__1
       (.I0(g0_b0_i_61__1_n_0),
        .I1(g0_b0_i_62__2_n_0),
        .O(g0_b0_i_25__1_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_25__2
       (.I0(g0_b0_i_61__2_n_0),
        .I1(g0_b0_i_62__4_n_0),
        .O(g0_b0_i_25__2_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_25__3
       (.I0(g0_b0_i_61__3_n_0),
        .I1(g0_b0_i_62__5_n_0),
        .O(g0_b0_i_25__3_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_25__4
       (.I0(g0_b0_i_61__4_n_0),
        .I1(g0_b0_i_62__6_n_0),
        .O(g0_b0_i_25__4_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_25__5
       (.I0(g0_b0_i_61__5_n_0),
        .I1(g0_b0_i_62__3_n_0),
        .O(g0_b0_i_25__5_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_25__6
       (.I0(g0_b0_i_61__6_n_0),
        .I1(g0_b0_i_62_n_0),
        .O(g0_b0_i_25__6_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_26
       (.I0(g0_b0_i_63_n_0),
        .I1(g0_b0_i_64_n_0),
        .O(g0_b0_i_26_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_26__0
       (.I0(g0_b0_i_63__0_n_0),
        .I1(g0_b0_i_64__0_n_0),
        .O(g0_b0_i_26__0_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_26__1
       (.I0(g0_b0_i_63__1_n_0),
        .I1(g0_b0_i_64__1_n_0),
        .O(g0_b0_i_26__1_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_26__2
       (.I0(g0_b0_i_63__2_n_0),
        .I1(g0_b0_i_64__2_n_0),
        .O(g0_b0_i_26__2_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_26__3
       (.I0(g0_b0_i_63__3_n_0),
        .I1(g0_b0_i_64__3_n_0),
        .O(g0_b0_i_26__3_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_26__4
       (.I0(g0_b0_i_63__4_n_0),
        .I1(g0_b0_i_64__4_n_0),
        .O(g0_b0_i_26__4_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_26__5
       (.I0(g0_b0_i_63__5_n_0),
        .I1(g0_b0_i_64__5_n_0),
        .O(g0_b0_i_26__5_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_26__6
       (.I0(g0_b0_i_63__6_n_0),
        .I1(g0_b0_i_64__6_n_0),
        .O(g0_b0_i_26__6_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_27
       (.I0(g0_b0_i_65__4_n_0),
        .I1(g0_b0_i_66__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_67__5_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_69__5_n_0),
        .O(g0_b0_i_27_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_27__0
       (.I0(g0_b0_i_124_n_0),
        .I1(g0_b0_i_79__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_80__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_78__6_n_0),
        .O(g0_b0_i_27__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_27__1
       (.I0(g0_b0_i_86__2_n_0),
        .I1(g0_b0_i_110__0_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_89__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_67__5_n_0),
        .O(g0_b0_i_27__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_27__2
       (.I0(\u1/p_14_in ),
        .I1(g0_b0_i_73__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_77__5_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_11_in ),
        .O(g0_b0_i_27__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_27__3
       (.I0(g0_b0_i_89__3_n_0),
        .I1(\u1/p_17_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_13_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(g0_b0_i_71__6_n_0),
        .O(g0_b0_i_27__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_27__4
       (.I0(\u1/p_17_in ),
        .I1(\u1/p_5_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_67__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_18_in ),
        .O(g0_b0_i_27__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_27__5
       (.I0(\u1/p_18_in ),
        .I1(\u1/p_2_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_5_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_19_in ),
        .O(g0_b0_i_27__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_27__6
       (.I0(g0_b0_i_102__2_n_0),
        .I1(g0_b0_i_65__4_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_87__3_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_72__6_n_0),
        .O(g0_b0_i_27__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_28
       (.I0(g0_b0_i_115_n_0),
        .I1(g0_b0_i_110__0_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_101__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_67__5_n_0),
        .O(g0_b0_i_28_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_28__0
       (.I0(g0_b0_i_70__6_n_0),
        .I1(g0_b0_i_71__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_72__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_73__6_n_0),
        .O(g0_b0_i_28__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_28__1
       (.I0(g0_b0_i_102__2_n_0),
        .I1(g0_b0_i_99__1_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_87__3_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_119_n_0),
        .O(g0_b0_i_28__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_28__2
       (.I0(\u1/p_7_in ),
        .I1(\u1/p_16_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_71__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_72__5_n_0),
        .O(g0_b0_i_28__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_28__3
       (.I0(\u1/p_9_in ),
        .I1(\u1/p_1_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_10_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(g0_b0_i_67__6_n_0),
        .O(g0_b0_i_28__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_28__4
       (.I0(g0_b0_i_98__1_n_0),
        .I1(\u1/p_15_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_0_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_96__2_n_0),
        .O(g0_b0_i_28__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_28__5
       (.I0(g0_b0_i_65__1_n_0),
        .I1(roundSel[0]),
        .I2(g0_b0_i_66__3_n_0),
        .I3(decrypt),
        .I4(g0_b0_i_67__4_n_0),
        .O(g0_b0_i_28__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_28__6
       (.I0(\u1/p_3_in ),
        .I1(\u1/p_7_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_74__6_n_0),
        .I4(g0_b0_i_75__6_n_0),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_28__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_29
       (.I0(g0_b0_i_80__6_n_0),
        .I1(g0_b0_i_99__1_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_77__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_119_n_0),
        .O(g0_b0_i_29_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_29__0
       (.I0(g0_b0_i_115_n_0),
        .I1(g0_b0_i_100__1_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_101__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_98__2_n_0),
        .O(g0_b0_i_29__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_29__1
       (.I0(g0_b0_i_66__5_n_0),
        .I1(g0_b0_i_72__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_73__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_70__6_n_0),
        .O(g0_b0_i_29__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_29__2
       (.I0(g0_b0_i_72__5_n_0),
        .I1(\u1/p_17_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_16_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(g0_b0_i_71__6_n_0),
        .O(g0_b0_i_29__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_29__3
       (.I0(g0_b0_i_73__5_n_0),
        .I1(g0_b0_i_74__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_75__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_3_in ),
        .O(g0_b0_i_29__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_29__4
       (.I0(\u1/p_14_in ),
        .I1(\u1/p_2_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_77__5_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_19_in ),
        .O(g0_b0_i_29__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_29__5
       (.I0(g0_b0_i_89__3_n_0),
        .I1(\u1/p_8_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_13_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_95__2_n_0),
        .O(g0_b0_i_29__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_29__6
       (.I0(g0_b0_i_74__5_n_0),
        .I1(roundSel[0]),
        .I2(g0_b0_i_75__5_n_0),
        .I3(decrypt),
        .I4(g0_b0_i_76__5_n_0),
        .O(g0_b0_i_29__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_2__0
       (.I0(desOut[17]),
        .I1(g0_b0_i_10__6_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_11__0_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_12__5_n_0),
        .O(\u0/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_2__1
       (.I0(desOut[51]),
        .I1(g0_b0_i_10__0_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_11__2_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_12__1_n_0),
        .O(\u0/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_2__2
       (.I0(desOut[19]),
        .I1(g0_b0_i_10__1_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_11__1_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_12__0_n_0),
        .O(\u0/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_2__3
       (.I0(desOut[53]),
        .I1(g0_b0_i_10__2_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_11__5_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_12__4_n_0),
        .O(\u0/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_2__4
       (.I0(desOut[55]),
        .I1(g0_b0_i_10__4_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_11__3_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_12__2_n_0),
        .O(\u0/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_2__5
       (.I0(desOut[21]),
        .I1(g0_b0_i_10__3_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_11__6_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_12__6_n_0),
        .O(\u0/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_2__6
       (.I0(desOut[23]),
        .I1(g0_b0_i_10__5_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_11__4_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_12__3_n_0),
        .O(\u0/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_3
       (.I0(desOut[41]),
        .I1(g0_b0_i_13_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_14_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_15_n_0),
        .O(\u0/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_30
       (.I0(g0_b0_i_77__6_n_0),
        .I1(g0_b0_i_78__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_79__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_80__6_n_0),
        .O(g0_b0_i_30_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_30__0
       (.I0(g0_b0_i_67__5_n_0),
        .I1(g0_b0_i_89__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_69__5_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_65__4_n_0),
        .O(g0_b0_i_30__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_30__1
       (.I0(g0_b0_i_78__6_n_0),
        .I1(g0_b0_i_80__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_77__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_90__3_n_0),
        .O(g0_b0_i_30__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_30__2
       (.I0(\u1/p_1_in ),
        .I1(\u1/p_18_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_5_in ),
        .I4(g0_b0_i_67__6_n_0),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_30__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_30__3
       (.I0(\u1/p_15_in ),
        .I1(\u1/p_3_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_74__6_n_0),
        .I4(g0_b0_i_96__2_n_0),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_30__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_30__4
       (.I0(g0_b0_i_77__5_n_0),
        .I1(\u1/p_8_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_11_in ),
        .I4(\u1/p_14_in ),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_30__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_30__5
       (.I0(g0_b0_i_73__5_n_0),
        .I1(\u1/p_9_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_10_in ),
        .I4(\u1/p_11_in ),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_30__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    g0_b0_i_30__6
       (.I0(g0_b0_i_65__2_n_0),
        .I1(decrypt),
        .I2(g0_b0_i_66__4_n_0),
        .I3(roundSel[0]),
        .I4(g0_b0_i_67__3_n_0),
        .O(g0_b0_i_30__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_31
       (.I0(g0_b0_i_68_n_0),
        .I1(g0_b0_i_69__0_n_0),
        .O(g0_b0_i_31_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_31__0
       (.I0(g0_b0_i_66_n_0),
        .I1(g0_b0_i_67_n_0),
        .O(g0_b0_i_31__0_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_31__1
       (.I0(g0_b0_i_68__0_n_0),
        .I1(g0_b0_i_69__1_n_0),
        .O(g0_b0_i_31__1_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_31__2
       (.I0(g0_b0_i_65_n_0),
        .I1(g0_b0_i_66__2_n_0),
        .O(g0_b0_i_31__2_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_31__3
       (.I0(g0_b0_i_81__0_n_0),
        .I1(g0_b0_i_82__2_n_0),
        .O(g0_b0_i_31__3_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_31__4
       (.I0(g0_b0_i_66__0_n_0),
        .I1(g0_b0_i_67__0_n_0),
        .O(g0_b0_i_31__4_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_31__5
       (.I0(g0_b0_i_65__0_n_0),
        .I1(g0_b0_i_66__1_n_0),
        .O(g0_b0_i_31__5_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_31__6
       (.I0(g0_b0_i_81__2_n_0),
        .I1(g0_b0_i_82__0_n_0),
        .O(g0_b0_i_31__6_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_32
       (.I0(g0_b0_i_83__0_n_0),
        .I1(g0_b0_i_84__0_n_0),
        .O(g0_b0_i_32_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_32__0
       (.I0(g0_b0_i_68__1_n_0),
        .I1(g0_b0_i_69__2_n_0),
        .O(g0_b0_i_32__0_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_32__1
       (.I0(g0_b0_i_70__2_n_0),
        .I1(g0_b0_i_71__3_n_0),
        .O(g0_b0_i_32__1_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_32__2
       (.I0(g0_b0_i_67__1_n_0),
        .I1(g0_b0_i_68__3_n_0),
        .O(g0_b0_i_32__2_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_32__3
       (.I0(g0_b0_i_83__1_n_0),
        .I1(g0_b0_i_84__1_n_0),
        .O(g0_b0_i_32__3_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_32__4
       (.I0(g0_b0_i_68__2_n_0),
        .I1(g0_b0_i_69__3_n_0),
        .O(g0_b0_i_32__4_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_32__5
       (.I0(g0_b0_i_67__2_n_0),
        .I1(g0_b0_i_68__4_n_0),
        .O(g0_b0_i_32__5_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_32__6
       (.I0(g0_b0_i_70__3_n_0),
        .I1(g0_b0_i_71__2_n_0),
        .O(g0_b0_i_32__6_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_33
       (.I0(g0_b0_i_67__5_n_0),
        .I1(g0_b0_i_73__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_110__0_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_66__5_n_0),
        .O(g0_b0_i_33_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_33__0
       (.I0(g0_b0_i_85__3_n_0),
        .I1(g0_b0_i_86__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_70__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_87__3_n_0),
        .O(g0_b0_i_33__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_33__1
       (.I0(g0_b0_i_69__5_n_0),
        .I1(g0_b0_i_99__1_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_66__5_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_119_n_0),
        .O(g0_b0_i_33__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    g0_b0_i_33__2
       (.I0(g0_b0_i_70__4_n_0),
        .I1(decrypt),
        .I2(g0_b0_i_71__4_n_0),
        .I3(roundSel[0]),
        .I4(g0_b0_i_72__0_n_0),
        .O(g0_b0_i_33__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_33__3
       (.I0(\u1/p_2_in ),
        .I1(g0_b0_i_74__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_96__2_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_3_in ),
        .O(g0_b0_i_33__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_33__4
       (.I0(g0_b0_i_71__6_n_0),
        .I1(\u1/p_18_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_17_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_0_in ),
        .O(g0_b0_i_33__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_33__5
       (.I0(g0_b0_i_75__6_n_0),
        .I1(g0_b0_i_98__1_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_7_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_13_in ),
        .O(g0_b0_i_33__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_33__6
       (.I0(\u1/p_19_in ),
        .I1(\u1/p_3_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_2_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_16_in ),
        .O(g0_b0_i_33__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    g0_b0_i_34
       (.I0(g0_b0_i_72__4_n_0),
        .I1(decrypt),
        .I2(g0_b0_i_73__4_n_0),
        .I3(roundSel[0]),
        .I4(g0_b0_i_74__4_n_0),
        .O(g0_b0_i_34_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_34__0
       (.I0(g0_b0_i_79__6_n_0),
        .I1(g0_b0_i_69__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_88__3_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_89__2_n_0),
        .O(g0_b0_i_34__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_34__1
       (.I0(g0_b0_i_73__6_n_0),
        .I1(g0_b0_i_88__3_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_71__5_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_79__6_n_0),
        .O(g0_b0_i_34__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_34__2
       (.I0(g0_b0_i_86__2_n_0),
        .I1(g0_b0_i_100__1_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_89__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_98__2_n_0),
        .O(g0_b0_i_34__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_34__3
       (.I0(\u1/p_11_in ),
        .I1(\u1/p_18_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_73__5_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_0_in ),
        .O(g0_b0_i_34__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_34__4
       (.I0(g0_b0_i_67__6_n_0),
        .I1(\u1/p_14_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_1_in ),
        .I4(g0_b0_i_74__6_n_0),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_34__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_34__5
       (.I0(\u1/p_1_in ),
        .I1(g0_b0_i_77__5_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_19_in ),
        .I4(\u1/p_14_in ),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_34__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_34__6
       (.I0(g0_b0_i_75__6_n_0),
        .I1(g0_b0_i_72__5_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_7_in ),
        .I4(\u1/p_5_in ),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_34__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_35
       (.I0(g0_b0_i_85__3_n_0),
        .I1(g0_b0_i_80__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_70__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_124_n_0),
        .O(g0_b0_i_35_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_35__0
       (.I0(g0_b0_i_90__3_n_0),
        .I1(g0_b0_i_73__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_78__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_66__5_n_0),
        .O(g0_b0_i_35__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_35__1
       (.I0(g0_b0_i_69__5_n_0),
        .I1(g0_b0_i_70__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_66__5_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_85__3_n_0),
        .O(g0_b0_i_35__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_35__2
       (.I0(g0_b0_i_102__2_n_0),
        .I1(g0_b0_i_78__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_87__3_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_90__3_n_0),
        .O(g0_b0_i_35__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_35__3
       (.I0(g0_b0_i_71__6_n_0),
        .I1(\u1/p_9_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_17_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_77__5_n_0),
        .O(g0_b0_i_35__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_35__4
       (.I0(\u1/p_17_in ),
        .I1(\u1/p_10_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_67__6_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_9_in ),
        .O(g0_b0_i_35__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_35__5
       (.I0(\u1/p_11_in ),
        .I1(\u1/p_3_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_73__5_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_16_in ),
        .O(g0_b0_i_35__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_35__6
       (.I0(g0_b0_i_95__2_n_0),
        .I1(g0_b0_i_72__5_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_8_in ),
        .I4(\u1/p_5_in ),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_35__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_36
       (.I0(g0_b0_i_115_n_0),
        .I1(g0_b0_i_79__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_88__3_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_77__6_n_0),
        .O(g0_b0_i_36_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_36__0
       (.I0(g0_b0_i_88__3_n_0),
        .I1(g0_b0_i_115_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_101__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_79__6_n_0),
        .O(g0_b0_i_36__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_36__1
       (.I0(g0_b0_i_65__4_n_0),
        .I1(g0_b0_i_86__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_89__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_72__6_n_0),
        .O(g0_b0_i_36__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_36__2
       (.I0(\u1/p_13_in ),
        .I1(\u1/p_7_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_71__6_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(g0_b0_i_89__3_n_0),
        .O(g0_b0_i_36__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_36__3
       (.I0(\u1/p_14_in ),
        .I1(g0_b0_i_95__2_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_8_in ),
        .I4(g0_b0_i_74__6_n_0),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_36__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_36__4
       (.I0(\u1/p_3_in ),
        .I1(g0_b0_i_96__2_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_15_in ),
        .I4(\u1/p_16_in ),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_36__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    g0_b0_i_36__5
       (.I0(g0_b0_i_91__3_n_0),
        .I1(decrypt),
        .I2(g0_b0_i_92__3_n_0),
        .I3(roundSel[0]),
        .I4(g0_b0_i_93__2_n_0),
        .O(g0_b0_i_36__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_36__6
       (.I0(g0_b0_i_89__3_n_0),
        .I1(g0_b0_i_75__6_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_7_in ),
        .I4(\u1/p_10_in ),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_36__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_37
       (.I0(g0_b0_i_75_n_0),
        .I1(g0_b0_i_76__0_n_0),
        .O(g0_b0_i_37_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_37__0
       (.I0(g0_b0_i_94_n_0),
        .I1(g0_b0_i_95_n_0),
        .O(g0_b0_i_37__0_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_37__1
       (.I0(g0_b0_i_73_n_0),
        .I1(g0_b0_i_74__0_n_0),
        .O(g0_b0_i_37__1_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_37__2
       (.I0(g0_b0_i_72_n_0),
        .I1(g0_b0_i_73__2_n_0),
        .O(g0_b0_i_37__2_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_37__3
       (.I0(g0_b0_i_69_n_0),
        .I1(g0_b0_i_70__0_n_0),
        .O(g0_b0_i_37__3_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_37__4
       (.I0(g0_b0_i_91__0_n_0),
        .I1(g0_b0_i_92__1_n_0),
        .O(g0_b0_i_37__4_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_37__5
       (.I0(g0_b0_i_70_n_0),
        .I1(g0_b0_i_71_n_0),
        .O(g0_b0_i_37__5_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_37__6
       (.I0(g0_b0_i_69__4_n_0),
        .I1(g0_b0_i_70__1_n_0),
        .O(g0_b0_i_37__6_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_38
       (.I0(g0_b0_i_77__2_n_0),
        .I1(g0_b0_i_78__3_n_0),
        .O(g0_b0_i_38_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_38__0
       (.I0(g0_b0_i_96__0_n_0),
        .I1(g0_b0_i_97_n_0),
        .O(g0_b0_i_38__0_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_38__1
       (.I0(g0_b0_i_75__1_n_0),
        .I1(g0_b0_i_76__2_n_0),
        .O(g0_b0_i_38__1_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_38__2
       (.I0(g0_b0_i_74__3_n_0),
        .I1(g0_b0_i_75__4_n_0),
        .O(g0_b0_i_38__2_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_38__3
       (.I0(g0_b0_i_72__1_n_0),
        .I1(g0_b0_i_73__3_n_0),
        .O(g0_b0_i_38__3_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_38__4
       (.I0(g0_b0_i_71__0_n_0),
        .I1(g0_b0_i_72__3_n_0),
        .O(g0_b0_i_38__4_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_38__5
       (.I0(g0_b0_i_71__1_n_0),
        .I1(g0_b0_i_72__2_n_0),
        .O(g0_b0_i_38__5_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_38__6
       (.I0(g0_b0_i_93__1_n_0),
        .I1(g0_b0_i_94__3_n_0),
        .O(g0_b0_i_38__6_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_39
       (.I0(g0_b0_i_78__6_n_0),
        .I1(g0_b0_i_101__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_79__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_115_n_0),
        .O(g0_b0_i_39_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_39__0
       (.I0(g0_b0_i_66__5_n_0),
        .I1(g0_b0_i_98__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_73__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_99__1_n_0),
        .O(g0_b0_i_39__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_39__1
       (.I0(g0_b0_i_87__3_n_0),
        .I1(g0_b0_i_67__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_86__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_65__4_n_0),
        .O(g0_b0_i_39__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_39__2
       (.I0(g0_b0_i_77__6_n_0),
        .I1(g0_b0_i_85__3_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_115_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_88__3_n_0),
        .O(g0_b0_i_39__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_39__3
       (.I0(\u1/p_0_in ),
        .I1(\u1/p_19_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_18_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_1_in ),
        .O(g0_b0_i_39__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_39__4
       (.I0(g0_b0_i_95__2_n_0),
        .I1(\u1/p_9_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_8_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_77__5_n_0),
        .O(g0_b0_i_39__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_39__5
       (.I0(g0_b0_i_77__5_n_0),
        .I1(g0_b0_i_75__6_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_9_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(g0_b0_i_73__5_n_0),
        .O(g0_b0_i_39__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_39__6
       (.I0(g0_b0_i_74__6_n_0),
        .I1(\u1/p_11_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_14_in ),
        .I4(\u1/p_8_in ),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_39__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_3__0
       (.I0(desOut[9]),
        .I1(g0_b0_i_13__0_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_14__0_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_15__0_n_0),
        .O(\u0/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_3__1
       (.I0(desOut[11]),
        .I1(g0_b0_i_13__2_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_14__1_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_15__1_n_0),
        .O(\u0/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_3__2
       (.I0(desOut[43]),
        .I1(g0_b0_i_13__1_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_14__2_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_15__2_n_0),
        .O(\u0/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_3__3
       (.I0(desOut[45]),
        .I1(g0_b0_i_13__3_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_14__3_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_15__3_n_0),
        .O(\u0/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_3__4
       (.I0(desOut[13]),
        .I1(g0_b0_i_13__4_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_14__4_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_15__4_n_0),
        .O(\u0/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_3__5
       (.I0(desOut[47]),
        .I1(g0_b0_i_13__5_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_14__5_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_15__5_n_0),
        .O(\u0/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_3__6
       (.I0(desOut[15]),
        .I1(g0_b0_i_13__6_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_14__6_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_15__6_n_0),
        .O(\u0/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_4
       (.I0(desOut[33]),
        .I1(g0_b0_i_16_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_17__6_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_18_n_0),
        .O(\u0/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_40
       (.I0(g0_b0_i_100__1_n_0),
        .I1(g0_b0_i_87__3_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_90__3_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_102__2_n_0),
        .O(g0_b0_i_40_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_40__0
       (.I0(g0_b0_i_89__2_n_0),
        .I1(g0_b0_i_90__3_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_69__5_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_100__1_n_0),
        .O(g0_b0_i_40__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_40__1
       (.I0(g0_b0_i_124_n_0),
        .I1(g0_b0_i_72__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_80__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_70__6_n_0),
        .O(g0_b0_i_40__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_40__2
       (.I0(g0_b0_i_101__2_n_0),
        .I1(g0_b0_i_119_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_102__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_110__0_n_0),
        .O(g0_b0_i_40__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_40__3
       (.I0(\u1/p_13_in ),
        .I1(g0_b0_i_96__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_98__1_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_2_in ),
        .O(g0_b0_i_40__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_40__4
       (.I0(g0_b0_i_96__2_n_0),
        .I1(g0_b0_i_89__3_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_15_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_10_in ),
        .O(g0_b0_i_40__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_40__5
       (.I0(\u1/p_16_in ),
        .I1(g0_b0_i_75__6_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_3_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_73__5_n_0),
        .O(g0_b0_i_40__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_40__6
       (.I0(g0_b0_i_74__6_n_0),
        .I1(g0_b0_i_71__6_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_14_in ),
        .I4(\u1/p_7_in ),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_40__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_41
       (.I0(g0_b0_i_99__1_n_0),
        .I1(g0_b0_i_89__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_98__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_86__2_n_0),
        .O(g0_b0_i_41_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_41__0
       (.I0(g0_b0_i_87__3_n_0),
        .I1(g0_b0_i_79__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_86__2_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_78__6_n_0),
        .O(g0_b0_i_41__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_41__1
       (.I0(g0_b0_i_77__6_n_0),
        .I1(g0_b0_i_98__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_115_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_99__1_n_0),
        .O(g0_b0_i_41__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_41__2
       (.I0(\u1/p_10_in ),
        .I1(g0_b0_i_95__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_89__3_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_15_in ),
        .O(g0_b0_i_41__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_41__3
       (.I0(\u1/p_19_in ),
        .I1(g0_b0_i_98__1_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_2_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_13_in ),
        .O(g0_b0_i_41__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_41__4
       (.I0(\u1/p_16_in ),
        .I1(g0_b0_i_67__6_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_3_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_17_in ),
        .O(g0_b0_i_41__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_41__5
       (.I0(\u1/p_5_in ),
        .I1(g0_b0_i_71__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_72__5_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_7_in ),
        .O(g0_b0_i_41__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_41__6
       (.I0(g0_b0_i_77__4_n_0),
        .I1(roundSel[0]),
        .I2(g0_b0_i_78__4_n_0),
        .I3(decrypt),
        .I4(g0_b0_i_79__4_n_0),
        .O(g0_b0_i_41__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_42
       (.I0(g0_b0_i_66__5_n_0),
        .I1(g0_b0_i_110__0_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_119_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_69__5_n_0),
        .O(g0_b0_i_42_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_42__0
       (.I0(g0_b0_i_85__3_n_0),
        .I1(g0_b0_i_101__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_102__2_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_88__3_n_0),
        .O(g0_b0_i_42__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_42__1
       (.I0(g0_b0_i_90__3_n_0),
        .I1(g0_b0_i_124_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_80__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_100__1_n_0),
        .O(g0_b0_i_42__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_42__2
       (.I0(g0_b0_i_119_n_0),
        .I1(g0_b0_i_66__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_73__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_110__0_n_0),
        .O(g0_b0_i_42__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_42__3
       (.I0(\u1/p_11_in ),
        .I1(g0_b0_i_77__5_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_9_in ),
        .I4(\u1/p_8_in ),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_42__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_42__4
       (.I0(\u1/p_18_in ),
        .I1(g0_b0_i_67__6_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_1_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_0_in ),
        .O(g0_b0_i_42__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_42__5
       (.I0(\u1/p_19_in ),
        .I1(\u1/p_5_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_72__5_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_1_in ),
        .O(g0_b0_i_42__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_42__6
       (.I0(g0_b0_i_67__6_n_0),
        .I1(\u1/p_0_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_18_in ),
        .I4(\u1/p_17_in ),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_42__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_43
       (.I0(g0_b0_i_79_n_0),
        .I1(g0_b0_i_80__1_n_0),
        .O(g0_b0_i_43_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_43__0
       (.I0(g0_b0_i_103_n_0),
        .I1(g0_b0_i_104_n_0),
        .O(g0_b0_i_43__0_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_43__1
       (.I0(g0_b0_i_80_n_0),
        .I1(g0_b0_i_81__3_n_0),
        .O(g0_b0_i_43__1_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_43__2
       (.I0(g0_b0_i_76_n_0),
        .I1(g0_b0_i_77__1_n_0),
        .O(g0_b0_i_43__2_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_43__3
       (.I0(g0_b0_i_73__0_n_0),
        .I1(g0_b0_i_74__2_n_0),
        .O(g0_b0_i_43__3_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_43__4
       (.I0(g0_b0_i_101_n_0),
        .I1(g0_b0_i_102_n_0),
        .O(g0_b0_i_43__4_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_43__5
       (.I0(g0_b0_i_74_n_0),
        .I1(g0_b0_i_75__0_n_0),
        .O(g0_b0_i_43__5_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_43__6
       (.I0(g0_b0_i_73__1_n_0),
        .I1(g0_b0_i_74__1_n_0),
        .O(g0_b0_i_43__6_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_44
       (.I0(g0_b0_i_81__5_n_0),
        .I1(g0_b0_i_82__5_n_0),
        .O(g0_b0_i_44_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_44__0
       (.I0(g0_b0_i_82__3_n_0),
        .I1(g0_b0_i_83__4_n_0),
        .O(g0_b0_i_44__0_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_44__1
       (.I0(g0_b0_i_78__2_n_0),
        .I1(g0_b0_i_79__3_n_0),
        .O(g0_b0_i_44__1_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_44__2
       (.I0(g0_b0_i_75__2_n_0),
        .I1(g0_b0_i_76__3_n_0),
        .O(g0_b0_i_44__2_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_44__3
       (.I0(g0_b0_i_103__0_n_0),
        .I1(g0_b0_i_104__0_n_0),
        .O(g0_b0_i_44__3_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_44__4
       (.I0(g0_b0_i_76__1_n_0),
        .I1(g0_b0_i_77__3_n_0),
        .O(g0_b0_i_44__4_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_44__5
       (.I0(g0_b0_i_75__3_n_0),
        .I1(g0_b0_i_76__4_n_0),
        .O(g0_b0_i_44__5_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_44__6
       (.I0(g0_b0_i_105__1_n_0),
        .I1(g0_b0_i_106__0_n_0),
        .O(g0_b0_i_44__6_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_45
       (.I0(\u1/p_16_in ),
        .I1(g0_b0_i_95__2_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_3_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_15_in ),
        .O(g0_b0_i_45_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_45__0
       (.I0(\u1/p_9_in ),
        .I1(\u1/p_7_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_10_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_75__6_n_0),
        .O(g0_b0_i_45__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_45__1
       (.I0(\u1/p_10_in ),
        .I1(g0_b0_i_71__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_89__3_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_7_in ),
        .O(g0_b0_i_45__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_45__2
       (.I0(g0_b0_i_67__6_n_0),
        .I1(g0_b0_i_72__5_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_1_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_5_in ),
        .O(g0_b0_i_45__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_45__3
       (.I0(g0_b0_i_80__6_n_0),
        .I1(g0_b0_i_88__3_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_77__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_79__6_n_0),
        .O(g0_b0_i_45__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    g0_b0_i_45__4
       (.I0(g0_b0_i_84__5_n_0),
        .I1(decrypt),
        .I2(g0_b0_i_85__1_n_0),
        .I3(roundSel[0]),
        .I4(g0_b0_i_86__0_n_0),
        .O(g0_b0_i_45__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_45__5
       (.I0(g0_b0_i_79__6_n_0),
        .I1(g0_b0_i_102__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_88__3_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_101__2_n_0),
        .O(g0_b0_i_45__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_45__6
       (.I0(g0_b0_i_83__5_n_0),
        .I1(roundSel[0]),
        .I2(g0_b0_i_92__3_n_0),
        .I3(decrypt),
        .I4(g0_b0_i_84__6_n_0),
        .O(g0_b0_i_45__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_46
       (.I0(g0_b0_i_110__0_n_0),
        .I1(g0_b0_i_77__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_119_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_80__6_n_0),
        .O(g0_b0_i_46_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    g0_b0_i_46__0
       (.I0(g0_b0_i_107__0_n_0),
        .I1(decrypt),
        .I2(g0_b0_i_108__0_n_0),
        .I3(roundSel[0]),
        .I4(g0_b0_i_109__0_n_0),
        .O(g0_b0_i_46__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_46__1
       (.I0(g0_b0_i_67__5_n_0),
        .I1(g0_b0_i_80__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_110__0_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_124_n_0),
        .O(g0_b0_i_46__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_46__2
       (.I0(g0_b0_i_90__3_n_0),
        .I1(g0_b0_i_86__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_78__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_87__3_n_0),
        .O(g0_b0_i_46__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_46__3
       (.I0(\u1/p_5_in ),
        .I1(\u1/p_11_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_72__5_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_8_in ),
        .O(g0_b0_i_46__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_46__4
       (.I0(g0_b0_i_77__5_n_0),
        .I1(g0_b0_i_67__6_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_9_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_17_in ),
        .O(g0_b0_i_46__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_46__5
       (.I0(g0_b0_i_71__6_n_0),
        .I1(\u1/p_3_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_17_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_16_in ),
        .O(g0_b0_i_46__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_46__6
       (.I0(\u1/p_14_in ),
        .I1(\u1/p_17_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_77__5_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_71__6_n_0),
        .O(g0_b0_i_46__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_47
       (.I0(g0_b0_i_65__4_n_0),
        .I1(g0_b0_i_101__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_67__5_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_115_n_0),
        .O(g0_b0_i_47_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_47__0
       (.I0(g0_b0_i_73__6_n_0),
        .I1(g0_b0_i_65__4_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_71__5_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_72__6_n_0),
        .O(g0_b0_i_47__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_47__1
       (.I0(g0_b0_i_72__6_n_0),
        .I1(g0_b0_i_115_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_65__4_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_77__6_n_0),
        .O(g0_b0_i_47__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_47__2
       (.I0(g0_b0_i_98__2_n_0),
        .I1(g0_b0_i_69__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_100__1_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_89__2_n_0),
        .O(g0_b0_i_47__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_47__3
       (.I0(\u1/p_0_in ),
        .I1(g0_b0_i_75__6_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_18_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(g0_b0_i_73__5_n_0),
        .O(g0_b0_i_47__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_47__4
       (.I0(g0_b0_i_74__6_n_0),
        .I1(\u1/p_19_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_14_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_1_in ),
        .O(g0_b0_i_47__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_47__5
       (.I0(g0_b0_i_75__6_n_0),
        .I1(\u1/p_14_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_7_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(g0_b0_i_74__6_n_0),
        .O(g0_b0_i_47__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_47__6
       (.I0(\u1/p_3_in ),
        .I1(\u1/p_1_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_74__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_67__6_n_0),
        .O(g0_b0_i_47__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_48
       (.I0(g0_b0_i_87__3_n_0),
        .I1(g0_b0_i_70__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_72__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_102__2_n_0),
        .O(g0_b0_i_48_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_48__0
       (.I0(g0_b0_i_71__6_n_0),
        .I1(\u1/p_13_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_98__1_n_0),
        .I4(\u1/p_7_in ),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_48__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_48__1
       (.I0(\u1/p_2_in ),
        .I1(g0_b0_i_72__5_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_16_in ),
        .I4(\u1/p_19_in ),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_48__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_48__2
       (.I0(g0_b0_i_96__2_n_0),
        .I1(\u1/p_16_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_3_in ),
        .I4(\u1/p_2_in ),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_48__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_48__3
       (.I0(\u1/p_9_in ),
        .I1(\u1/p_11_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_73__5_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(g0_b0_i_77__5_n_0),
        .O(g0_b0_i_48__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_48__4
       (.I0(g0_b0_i_110__0_n_0),
        .I1(g0_b0_i_69__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_66__5_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_67__5_n_0),
        .O(g0_b0_i_48__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_48__5
       (.I0(g0_b0_i_102__2_n_0),
        .I1(g0_b0_i_85__3_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_70__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_101__2_n_0),
        .O(g0_b0_i_48__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_48__6
       (.I0(g0_b0_i_73__6_n_0),
        .I1(g0_b0_i_119_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_99__1_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_66__5_n_0),
        .O(g0_b0_i_48__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_49
       (.I0(g0_b0_i_85_n_0),
        .I1(g0_b0_i_86_n_0),
        .O(g0_b0_i_49_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_49__0
       (.I0(g0_b0_i_111_n_0),
        .I1(g0_b0_i_112_n_0),
        .O(g0_b0_i_49__0_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_49__1
       (.I0(g0_b0_i_87_n_0),
        .I1(g0_b0_i_88_n_0),
        .O(g0_b0_i_49__1_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_49__2
       (.I0(g0_b0_i_80__0_n_0),
        .I1(g0_b0_i_81__4_n_0),
        .O(g0_b0_i_49__2_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_49__3
       (.I0(g0_b0_i_77_n_0),
        .I1(g0_b0_i_78__0_n_0),
        .O(g0_b0_i_49__3_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_49__4
       (.I0(g0_b0_i_105__0_n_0),
        .I1(g0_b0_i_106_n_0),
        .O(g0_b0_i_49__4_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_49__5
       (.I0(g0_b0_i_78_n_0),
        .I1(g0_b0_i_79__0_n_0),
        .O(g0_b0_i_49__5_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_49__6
       (.I0(g0_b0_i_77__0_n_0),
        .I1(g0_b0_i_78__1_n_0),
        .O(g0_b0_i_49__6_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_4__0
       (.I0(desOut[1]),
        .I1(g0_b0_i_16__0_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_17__3_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_18__4_n_0),
        .O(\u0/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_4__1
       (.I0(desOut[35]),
        .I1(g0_b0_i_16__1_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_17__4_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_18__5_n_0),
        .O(\u0/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_4__2
       (.I0(desOut[3]),
        .I1(g0_b0_i_16__2_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_17__5_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_18__6_n_0),
        .O(\u0/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_4__3
       (.I0(desOut[37]),
        .I1(g0_b0_i_16__3_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_17_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_18__0_n_0),
        .O(\u0/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_4__4
       (.I0(desOut[5]),
        .I1(g0_b0_i_16__4_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_17__1_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_18__2_n_0),
        .O(\u0/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_4__5
       (.I0(desOut[39]),
        .I1(g0_b0_i_16__5_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_17__2_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_18__3_n_0),
        .O(\u0/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_4__6
       (.I0(desOut[7]),
        .I1(g0_b0_i_16__6_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_17__0_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_18__1_n_0),
        .O(\u0/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_5
       (.I0(desOut[7]),
        .I1(g0_b0_i_19_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_20_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_21_n_0),
        .O(\u0/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_50
       (.I0(g0_b0_i_87__1_n_0),
        .I1(g0_b0_i_88__1_n_0),
        .O(g0_b0_i_50_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_50__0
       (.I0(g0_b0_i_113_n_0),
        .I1(g0_b0_i_114_n_0),
        .O(g0_b0_i_50__0_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_50__1
       (.I0(g0_b0_i_89_n_0),
        .I1(g0_b0_i_90_n_0),
        .O(g0_b0_i_50__1_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_50__2
       (.I0(g0_b0_i_82__4_n_0),
        .I1(g0_b0_i_83__3_n_0),
        .O(g0_b0_i_50__2_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_50__3
       (.I0(g0_b0_i_79__1_n_0),
        .I1(g0_b0_i_80__3_n_0),
        .O(g0_b0_i_50__3_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_50__4
       (.I0(g0_b0_i_107_n_0),
        .I1(g0_b0_i_108_n_0),
        .O(g0_b0_i_50__4_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_50__5
       (.I0(g0_b0_i_80__2_n_0),
        .I1(g0_b0_i_81__6_n_0),
        .O(g0_b0_i_50__5_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_50__6
       (.I0(g0_b0_i_79__2_n_0),
        .I1(g0_b0_i_80__4_n_0),
        .O(g0_b0_i_50__6_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_51
       (.I0(g0_b0_i_72__6_n_0),
        .I1(g0_b0_i_69__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_65__4_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_89__2_n_0),
        .O(g0_b0_i_51_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_51__0
       (.I0(g0_b0_i_90__3_n_0),
        .I1(g0_b0_i_115_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_78__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_77__6_n_0),
        .O(g0_b0_i_51__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_51__1
       (.I0(g0_b0_i_115_n_0),
        .I1(g0_b0_i_70__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_101__2_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_85__3_n_0),
        .O(g0_b0_i_51__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_51__2
       (.I0(g0_b0_i_101__2_n_0),
        .I1(g0_b0_i_72__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_102__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_70__6_n_0),
        .O(g0_b0_i_51__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_51__3
       (.I0(\u1/p_1_in ),
        .I1(\u1/p_16_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_19_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(g0_b0_i_72__5_n_0),
        .O(g0_b0_i_51__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_51__4
       (.I0(g0_b0_i_72__5_n_0),
        .I1(\u1/p_15_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_16_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_96__2_n_0),
        .O(g0_b0_i_51__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_51__5
       (.I0(\u1/p_15_in ),
        .I1(g0_b0_i_77__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_95__2_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_14_in ),
        .O(g0_b0_i_51__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_51__6
       (.I0(g0_b0_i_96__2_n_0),
        .I1(\u1/p_14_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_15_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_74__6_n_0),
        .O(g0_b0_i_51__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_52
       (.I0(g0_b0_i_85__3_n_0),
        .I1(g0_b0_i_73__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_70__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_66__5_n_0),
        .O(g0_b0_i_52_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_52__0
       (.I0(g0_b0_i_80__6_n_0),
        .I1(g0_b0_i_65__4_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_77__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_72__6_n_0),
        .O(g0_b0_i_52__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_52__1
       (.I0(g0_b0_i_98__2_n_0),
        .I1(g0_b0_i_102__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_100__1_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_101__2_n_0),
        .O(g0_b0_i_52__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_52__2
       (.I0(g0_b0_i_77__6_n_0),
        .I1(g0_b0_i_67__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_115_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_65__4_n_0),
        .O(g0_b0_i_52__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_52__3
       (.I0(\u1/p_17_in ),
        .I1(g0_b0_i_74__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_67__6_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_3_in ),
        .O(g0_b0_i_52__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_52__4
       (.I0(\u1/p_19_in ),
        .I1(\u1/p_9_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_2_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_77__5_n_0),
        .O(g0_b0_i_52__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_52__5
       (.I0(\u1/p_2_in ),
        .I1(\u1/p_10_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_96__2_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_9_in ),
        .O(g0_b0_i_52__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_52__6
       (.I0(\u1/p_18_in ),
        .I1(\u1/p_8_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_5_in ),
        .I4(g0_b0_i_95__2_n_0),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_52__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    g0_b0_i_53
       (.I0(g0_b0_i_89__1_n_0),
        .I1(decrypt),
        .I2(g0_b0_i_90__1_n_0),
        .I3(roundSel[0]),
        .I4(g0_b0_i_91__1_n_0),
        .O(g0_b0_i_53_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    g0_b0_i_53__0
       (.I0(g0_b0_i_116_n_0),
        .I1(decrypt),
        .I2(g0_b0_i_117_n_0),
        .I3(roundSel[0]),
        .I4(g0_b0_i_118_n_0),
        .O(g0_b0_i_53__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_53__1
       (.I0(g0_b0_i_119_n_0),
        .I1(g0_b0_i_86__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_99__1_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_87__3_n_0),
        .O(g0_b0_i_53__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_53__2
       (.I0(g0_b0_i_124_n_0),
        .I1(g0_b0_i_119_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_80__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_110__0_n_0),
        .O(g0_b0_i_53__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_53__3
       (.I0(\u1/p_7_in ),
        .I1(g0_b0_i_77__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_71__6_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_14_in ),
        .O(g0_b0_i_53__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_53__4
       (.I0(g0_b0_i_67__6_n_0),
        .I1(g0_b0_i_89__3_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_1_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_10_in ),
        .O(g0_b0_i_53__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_53__5
       (.I0(\u1/p_1_in ),
        .I1(\u1/p_13_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_19_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(g0_b0_i_89__3_n_0),
        .O(g0_b0_i_53__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_53__6
       (.I0(g0_b0_i_98__1_n_0),
        .I1(g0_b0_i_73__5_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_0_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_11_in ),
        .O(g0_b0_i_53__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_54
       (.I0(g0_b0_i_80__6_n_0),
        .I1(g0_b0_i_90__3_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_78__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_124_n_0),
        .O(g0_b0_i_54_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_54__0
       (.I0(g0_b0_i_69__5_n_0),
        .I1(g0_b0_i_67__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_110__0_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_89__2_n_0),
        .O(g0_b0_i_54__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_54__1
       (.I0(g0_b0_i_99__1_n_0),
        .I1(g0_b0_i_73__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_71__5_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_119_n_0),
        .O(g0_b0_i_54__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_54__2
       (.I0(g0_b0_i_84__2_n_0),
        .I1(roundSel[0]),
        .I2(g0_b0_i_85__2_n_0),
        .I3(decrypt),
        .I4(g0_b0_i_86__1_n_0),
        .O(g0_b0_i_54__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_54__3
       (.I0(\u1/p_10_in ),
        .I1(g0_b0_i_73__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_75__6_n_0),
        .I4(\u1/p_9_in ),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_54__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_54__4
       (.I0(\u1/p_7_in ),
        .I1(g0_b0_i_89__3_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_13_in ),
        .I4(g0_b0_i_75__6_n_0),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_54__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_54__5
       (.I0(\u1/p_0_in ),
        .I1(\u1/p_17_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_67__6_n_0),
        .I4(g0_b0_i_98__1_n_0),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_54__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_54__6
       (.I0(g0_b0_i_98__1_n_0),
        .I1(g0_b0_i_71__6_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_17_in ),
        .I4(\u1/p_13_in ),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_54__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_55
       (.I0(g0_b0_i_92_n_0),
        .I1(g0_b0_i_93_n_0),
        .O(g0_b0_i_55_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_55__0
       (.I0(g0_b0_i_120_n_0),
        .I1(g0_b0_i_121_n_0),
        .O(g0_b0_i_55__0_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_55__1
       (.I0(g0_b0_i_91_n_0),
        .I1(g0_b0_i_92__0_n_0),
        .O(g0_b0_i_55__1_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_55__2
       (.I0(g0_b0_i_87__0_n_0),
        .I1(g0_b0_i_88__0_n_0),
        .O(g0_b0_i_55__2_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_55__3
       (.I0(g0_b0_i_81_n_0),
        .I1(g0_b0_i_82__1_n_0),
        .O(g0_b0_i_55__3_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_55__4
       (.I0(g0_b0_i_109_n_0),
        .I1(g0_b0_i_110_n_0),
        .O(g0_b0_i_55__4_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_55__5
       (.I0(g0_b0_i_82_n_0),
        .I1(g0_b0_i_83_n_0),
        .O(g0_b0_i_55__5_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_55__6
       (.I0(g0_b0_i_81__1_n_0),
        .I1(g0_b0_i_82__6_n_0),
        .O(g0_b0_i_55__6_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_56
       (.I0(g0_b0_i_94__1_n_0),
        .I1(g0_b0_i_95__0_n_0),
        .O(g0_b0_i_56_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_56__0
       (.I0(g0_b0_i_122_n_0),
        .I1(g0_b0_i_123_n_0),
        .O(g0_b0_i_56__0_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_56__1
       (.I0(g0_b0_i_93__0_n_0),
        .I1(g0_b0_i_94__2_n_0),
        .O(g0_b0_i_56__1_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_56__2
       (.I0(g0_b0_i_89__0_n_0),
        .I1(g0_b0_i_90__0_n_0),
        .O(g0_b0_i_56__2_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_56__3
       (.I0(g0_b0_i_111__0_n_0),
        .I1(g0_b0_i_112__0_n_0),
        .O(g0_b0_i_56__3_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_56__4
       (.I0(g0_b0_i_83__2_n_0),
        .I1(g0_b0_i_84__3_n_0),
        .O(g0_b0_i_56__4_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_56__5
       (.I0(g0_b0_i_84_n_0),
        .I1(g0_b0_i_85__0_n_0),
        .O(g0_b0_i_56__5_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_56__6
       (.I0(g0_b0_i_83__6_n_0),
        .I1(g0_b0_i_84__4_n_0),
        .O(g0_b0_i_56__6_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_57
       (.I0(g0_b0_i_100__1_n_0),
        .I1(g0_b0_i_77__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_90__3_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_80__6_n_0),
        .O(g0_b0_i_57_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_57__0
       (.I0(g0_b0_i_70__6_n_0),
        .I1(g0_b0_i_89__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_72__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_86__2_n_0),
        .O(g0_b0_i_57__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_57__1
       (.I0(g0_b0_i_98__2_n_0),
        .I1(g0_b0_i_80__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_100__1_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_124_n_0),
        .O(g0_b0_i_57__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_57__2
       (.I0(g0_b0_i_73__6_n_0),
        .I1(g0_b0_i_100__1_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_71__5_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_98__2_n_0),
        .O(g0_b0_i_57__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_57__3
       (.I0(\u1/p_11_in ),
        .I1(g0_b0_i_89__3_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_73__5_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_10_in ),
        .O(g0_b0_i_57__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_57__4
       (.I0(\u1/p_8_in ),
        .I1(\u1/p_10_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_11_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_9_in ),
        .O(g0_b0_i_57__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_57__5
       (.I0(\u1/p_5_in ),
        .I1(g0_b0_i_96__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_72__5_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_2_in ),
        .O(g0_b0_i_57__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_57__6
       (.I0(\u1/p_13_in ),
        .I1(g0_b0_i_67__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_98__1_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_17_in ),
        .O(g0_b0_i_57__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_58
       (.I0(g0_b0_i_99__1_n_0),
        .I1(g0_b0_i_101__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_98__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_115_n_0),
        .O(g0_b0_i_58_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_58__0
       (.I0(g0_b0_i_119_n_0),
        .I1(g0_b0_i_115_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_99__1_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_77__6_n_0),
        .O(g0_b0_i_58__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_58__1
       (.I0(g0_b0_i_88__3_n_0),
        .I1(g0_b0_i_66__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_85__3_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_69__5_n_0),
        .O(g0_b0_i_58__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_58__2
       (.I0(g0_b0_i_69__5_n_0),
        .I1(g0_b0_i_78__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_66__5_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_90__3_n_0),
        .O(g0_b0_i_58__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_58__3
       (.I0(g0_b0_i_95__2_n_0),
        .I1(g0_b0_i_98__1_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_8_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_13_in ),
        .O(g0_b0_i_58__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_58__4
       (.I0(\u1/p_0_in ),
        .I1(g0_b0_i_95__2_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_18_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_15_in ),
        .O(g0_b0_i_58__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_58__5
       (.I0(\u1/p_10_in ),
        .I1(\u1/p_19_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_89__3_n_0),
        .I4(\u1/p_1_in ),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_58__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_58__6
       (.I0(\u1/p_15_in ),
        .I1(\u1/p_13_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_95__2_n_0),
        .I4(g0_b0_i_89__3_n_0),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_58__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_59
       (.I0(g0_b0_i_110__0_n_0),
        .I1(g0_b0_i_87__3_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_119_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_102__2_n_0),
        .O(g0_b0_i_59_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_59__0
       (.I0(g0_b0_i_67__5_n_0),
        .I1(g0_b0_i_102__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_110__0_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_101__2_n_0),
        .O(g0_b0_i_59__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_59__1
       (.I0(g0_b0_i_78__6_n_0),
        .I1(g0_b0_i_71__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_79__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_73__6_n_0),
        .O(g0_b0_i_59__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_59__2
       (.I0(g0_b0_i_86__2_n_0),
        .I1(g0_b0_i_88__3_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_89__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_79__6_n_0),
        .O(g0_b0_i_59__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_59__3
       (.I0(g0_b0_i_96__2_n_0),
        .I1(\u1/p_18_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_15_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_0_in ),
        .O(g0_b0_i_59__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_59__4
       (.I0(g0_b0_i_77__5_n_0),
        .I1(g0_b0_i_96__2_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_9_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_2_in ),
        .O(g0_b0_i_59__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_59__5
       (.I0(\u1/p_13_in ),
        .I1(\u1/p_11_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_98__1_n_0),
        .I4(\u1/p_8_in ),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_59__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_59__6
       (.I0(\u1/p_2_in ),
        .I1(\u1/p_0_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_96__2_n_0),
        .I4(g0_b0_i_98__1_n_0),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_59__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_5__0
       (.I0(desOut[33]),
        .I1(g0_b0_i_19__0_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_20__1_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_21__1_n_0),
        .O(\u0/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_5__1
       (.I0(desOut[1]),
        .I1(g0_b0_i_19__1_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_20__0_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_21__0_n_0),
        .O(\u0/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_5__2
       (.I0(desOut[35]),
        .I1(g0_b0_i_19__2_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_20__2_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_21__2_n_0),
        .O(\u0/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_5__3
       (.I0(desOut[3]),
        .I1(g0_b0_i_19__3_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_20__3_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_21__3_n_0),
        .O(\u0/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_5__4
       (.I0(desOut[37]),
        .I1(g0_b0_i_19__4_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_20__6_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_21__6_n_0),
        .O(\u0/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_5__5
       (.I0(desOut[39]),
        .I1(g0_b0_i_19__6_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_20__4_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_21__4_n_0),
        .O(\u0/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_5__6
       (.I0(desOut[5]),
        .I1(g0_b0_i_19__5_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_20__5_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_21__5_n_0),
        .O(\u0/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_6
       (.I0(desOut[25]),
        .I1(g0_b0_i_22_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_23_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_24_n_0),
        .O(\u0/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_60
       (.I0(g0_b0_i_89__2_n_0),
        .I1(g0_b0_i_65__4_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_67__5_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_86__2_n_0),
        .O(g0_b0_i_60_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_60__0
       (.I0(g0_b0_i_95__1_n_0),
        .I1(roundSel[0]),
        .I2(g0_b0_i_96__1_n_0),
        .I3(decrypt),
        .I4(g0_b0_i_97__1_n_0),
        .O(g0_b0_i_60__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_60__1
       (.I0(g0_b0_i_86__2_n_0),
        .I1(g0_b0_i_72__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_65__4_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_87__3_n_0),
        .O(g0_b0_i_60__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_60__2
       (.I0(g0_b0_i_70__6_n_0),
        .I1(g0_b0_i_102__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_87__3_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_85__3_n_0),
        .O(g0_b0_i_60__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_60__3
       (.I0(g0_b0_i_72__5_n_0),
        .I1(\u1/p_19_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_2_in ),
        .I4(\u1/p_5_in ),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_60__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_60__4
       (.I0(\u1/p_5_in ),
        .I1(\u1/p_1_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_19_in ),
        .I4(\u1/p_18_in ),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_60__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_60__5
       (.I0(g0_b0_i_75__6_n_0),
        .I1(\u1/p_10_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_89__3_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(g0_b0_i_73__5_n_0),
        .O(g0_b0_i_60__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_60__6
       (.I0(g0_b0_i_95__2_n_0),
        .I1(g0_b0_i_74__6_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_14_in ),
        .I4(\u1/p_15_in ),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_60__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_61
       (.I0(g0_b0_i_80__6_n_0),
        .I1(g0_b0_i_79__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_78__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_77__6_n_0),
        .O(g0_b0_i_61_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_61__0
       (.I0(g0_b0_i_90__3_n_0),
        .I1(g0_b0_i_77__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_80__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_78__6_n_0),
        .O(g0_b0_i_61__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_61__1
       (.I0(g0_b0_i_65__4_n_0),
        .I1(g0_b0_i_69__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_89__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_67__5_n_0),
        .O(g0_b0_i_61__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_61__2
       (.I0(g0_b0_i_67__6_n_0),
        .I1(\u1/p_5_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_18_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_1_in ),
        .O(g0_b0_i_61__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_61__3
       (.I0(\u1/p_14_in ),
        .I1(\u1/p_11_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_8_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_77__5_n_0),
        .O(g0_b0_i_61__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_61__4
       (.I0(g0_b0_i_96__2_n_0),
        .I1(g0_b0_i_74__6_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_3_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_15_in ),
        .O(g0_b0_i_61__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_61__5
       (.I0(\u1/p_11_in ),
        .I1(\u1/p_10_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_9_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_73__5_n_0),
        .O(g0_b0_i_61__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_61__6
       (.I0(g0_b0_i_96_n_0),
        .I1(roundSel[0]),
        .I2(g0_b0_i_97__0_n_0),
        .I3(decrypt),
        .I4(g0_b0_i_65__2_n_0),
        .O(g0_b0_i_61__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_62
       (.I0(g0_b0_i_119_n_0),
        .I1(g0_b0_i_77__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_99__1_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_80__6_n_0),
        .O(g0_b0_i_62_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    g0_b0_i_62__0
       (.I0(g0_b0_i_125_n_0),
        .I1(decrypt),
        .I2(g0_b0_i_75__5_n_0),
        .I3(roundSel[0]),
        .I4(g0_b0_i_126_n_0),
        .O(g0_b0_i_62__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_62__1
       (.I0(g0_b0_i_98__2_n_0),
        .I1(g0_b0_i_101__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_100__1_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_115_n_0),
        .O(g0_b0_i_62__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_62__2
       (.I0(g0_b0_i_70__6_n_0),
        .I1(g0_b0_i_73__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_72__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_66__5_n_0),
        .O(g0_b0_i_62__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_62__3
       (.I0(g0_b0_i_95__2_n_0),
        .I1(\u1/p_13_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_8_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_89__3_n_0),
        .O(g0_b0_i_62__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_62__4
       (.I0(g0_b0_i_71__6_n_0),
        .I1(\u1/p_16_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_17_in ),
        .I4(g0_b0_i_72__5_n_0),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_62__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_62__5
       (.I0(\u1/p_3_in ),
        .I1(g0_b0_i_75__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_74__6_n_0),
        .I4(g0_b0_i_73__5_n_0),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_62__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_62__6
       (.I0(\u1/p_19_in ),
        .I1(g0_b0_i_77__5_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_2_in ),
        .I4(\u1/p_14_in ),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_62__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_63
       (.I0(g0_b0_i_67__5_n_0),
        .I1(g0_b0_i_101__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_110__0_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_115_n_0),
        .O(g0_b0_i_63_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_63__0
       (.I0(g0_b0_i_73__6_n_0),
        .I1(g0_b0_i_72__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_71__5_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_70__6_n_0),
        .O(g0_b0_i_63__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_63__1
       (.I0(g0_b0_i_119_n_0),
        .I1(g0_b0_i_87__3_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_99__1_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_102__2_n_0),
        .O(g0_b0_i_63__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    g0_b0_i_63__2
       (.I0(g0_b0_i_67__4_n_0),
        .I1(decrypt),
        .I2(g0_b0_i_91__2_n_0),
        .I3(roundSel[0]),
        .I4(g0_b0_i_92__2_n_0),
        .O(g0_b0_i_63__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_63__3
       (.I0(g0_b0_i_75__6_n_0),
        .I1(g0_b0_i_74__6_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_7_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_3_in ),
        .O(g0_b0_i_63__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_63__4
       (.I0(g0_b0_i_72__5_n_0),
        .I1(g0_b0_i_71__6_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_16_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_7_in ),
        .O(g0_b0_i_63__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_63__5
       (.I0(g0_b0_i_67__6_n_0),
        .I1(\u1/p_10_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_1_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_9_in ),
        .O(g0_b0_i_63__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_63__6
       (.I0(g0_b0_i_96__2_n_0),
        .I1(\u1/p_0_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_15_in ),
        .I4(g0_b0_i_98__1_n_0),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_63__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_64
       (.I0(g0_b0_i_72__6_n_0),
        .I1(g0_b0_i_87__3_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_65__4_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_102__2_n_0),
        .O(g0_b0_i_64_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_64__0
       (.I0(g0_b0_i_69__5_n_0),
        .I1(g0_b0_i_67__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_66__5_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_65__4_n_0),
        .O(g0_b0_i_64__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_64__1
       (.I0(g0_b0_i_67__5_n_0),
        .I1(g0_b0_i_89__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_110__0_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_86__2_n_0),
        .O(g0_b0_i_64__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_64__2
       (.I0(g0_b0_i_78__6_n_0),
        .I1(g0_b0_i_80__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_79__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_124_n_0),
        .O(g0_b0_i_64__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_64__3
       (.I0(\u1/p_11_in ),
        .I1(g0_b0_i_77__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_73__5_n_0),
        .I4(\u1/p_14_in ),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_64__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_64__4
       (.I0(\u1/p_18_in ),
        .I1(g0_b0_i_67__6_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_5_in ),
        .I4(\u1/p_17_in ),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_64__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_64__5
       (.I0(g0_b0_i_71__6_n_0),
        .I1(\u1/p_13_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_17_in ),
        .I4(g0_b0_i_89__3_n_0),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_64__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_64__6
       (.I0(\u1/p_19_in ),
        .I1(\u1/p_5_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_2_in ),
        .I4(\u1/p_18_in ),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_64__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_65
       (.I0(\u1/p_16_in ),
        .I1(\u1/p_15_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_96__2_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_3_in ),
        .O(g0_b0_i_65_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_65__0
       (.I0(g0_b0_i_74__6_n_0),
        .I1(\u1/p_8_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_95__2_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_14_in ),
        .O(g0_b0_i_65__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_65__1
       (.I0(g0_b0_i_71__5_n_0),
        .I1(\u1/decrypt_int__2 ),
        .I2(g0_b0_i_85__3_n_0),
        .O(g0_b0_i_65__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFB08)) 
    g0_b0_i_65__2
       (.I0(key2[0]),
        .I1(roundSel[4]),
        .I2(roundSel[5]),
        .I3(g0_b0_i_100__1_n_0),
        .O(g0_b0_i_65__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB4)) 
    g0_b0_i_65__3
       (.I0(roundSel[5]),
        .I1(roundSel[4]),
        .I2(decrypt),
        .O(\u1/decrypt_int__2 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_65__4
       (.I0(key2[9]),
        .I1(roundSel[5]),
        .I2(key3[9]),
        .I3(decrypt),
        .I4(key1[9]),
        .I5(roundSel[4]),
        .O(g0_b0_i_65__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_65__5
       (.I0(key2[12]),
        .I1(roundSel[5]),
        .I2(key3[12]),
        .I3(decrypt),
        .I4(key1[12]),
        .I5(roundSel[4]),
        .O(\u1/p_17_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB4)) 
    g0_b0_i_65__6
       (.I0(roundSel[5]),
        .I1(roundSel[4]),
        .I2(decrypt),
        .O(g0_b0_i_65__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_66
       (.I0(g0_b0_i_72__6_n_0),
        .I1(g0_b0_i_89__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_86__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_65__4_n_0),
        .O(g0_b0_i_66_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_66__0
       (.I0(g0_b0_i_89__3_n_0),
        .I1(g0_b0_i_71__6_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_7_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_13_in ),
        .O(g0_b0_i_66__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_66__1
       (.I0(\u1/p_16_in ),
        .I1(g0_b0_i_73__5_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_3_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_11_in ),
        .O(g0_b0_i_66__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_66__2
       (.I0(\u1/p_5_in ),
        .I1(\u1/p_8_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_72__5_n_0),
        .I4(g0_b0_i_95__2_n_0),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_66__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_66__3
       (.I0(key1[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_88__3_n_0),
        .I3(roundSel[4]),
        .I4(key3[0]),
        .O(g0_b0_i_66__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_66__4
       (.I0(key3[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_100__1_n_0),
        .I3(roundSel[4]),
        .I4(key1[0]),
        .O(g0_b0_i_66__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_66__5
       (.I0(key2[44]),
        .I1(roundSel[5]),
        .I2(key3[44]),
        .I3(decrypt),
        .I4(key1[44]),
        .I5(roundSel[4]),
        .O(g0_b0_i_66__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_66__6
       (.I0(key2[47]),
        .I1(roundSel[5]),
        .I2(key3[47]),
        .I3(decrypt),
        .I4(key1[47]),
        .I5(roundSel[4]),
        .O(\u1/p_5_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_67
       (.I0(g0_b0_i_85__3_n_0),
        .I1(g0_b0_i_66__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_70__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_69__5_n_0),
        .O(g0_b0_i_67_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_67__0
       (.I0(\u1/p_9_in ),
        .I1(g0_b0_i_67__6_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_10_in ),
        .I4(\u1/p_17_in ),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_67__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_67__1
       (.I0(\u1/p_0_in ),
        .I1(g0_b0_i_73__5_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_18_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_11_in ),
        .O(g0_b0_i_67__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_67__2
       (.I0(\u1/p_5_in ),
        .I1(\u1/p_7_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_72__5_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_75__6_n_0),
        .O(g0_b0_i_67__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_67__3
       (.I0(g0_b0_i_124_n_0),
        .I1(\u1/decrypt_int__2 ),
        .I2(g0_b0_i_98__2_n_0),
        .O(g0_b0_i_67__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFB08)) 
    g0_b0_i_67__4
       (.I0(key2[0]),
        .I1(roundSel[4]),
        .I2(roundSel[5]),
        .I3(g0_b0_i_88__3_n_0),
        .O(g0_b0_i_67__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_67__5
       (.I0(key2[23]),
        .I1(roundSel[5]),
        .I2(key3[23]),
        .I3(decrypt),
        .I4(key1[23]),
        .I5(roundSel[4]),
        .O(g0_b0_i_67__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_67__6
       (.I0(key2[26]),
        .I1(roundSel[5]),
        .I2(key3[26]),
        .I3(decrypt),
        .I4(key1[26]),
        .I5(roundSel[4]),
        .O(g0_b0_i_67__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_68
       (.I0(g0_b0_i_77__6_n_0),
        .I1(g0_b0_i_88__3_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_79__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_115_n_0),
        .O(g0_b0_i_68_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_68__0
       (.I0(g0_b0_i_79__6_n_0),
        .I1(g0_b0_i_101__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_115_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_88__3_n_0),
        .O(g0_b0_i_68__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_68__1
       (.I0(g0_b0_i_79__6_n_0),
        .I1(g0_b0_i_71__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_88__3_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_73__6_n_0),
        .O(g0_b0_i_68__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_68__2
       (.I0(\u1/p_14_in ),
        .I1(\u1/p_19_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_77__5_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_1_in ),
        .O(g0_b0_i_68__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_68__3
       (.I0(\u1/p_13_in ),
        .I1(\u1/p_7_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_98__1_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(g0_b0_i_75__6_n_0),
        .O(g0_b0_i_68__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_68__4
       (.I0(\u1/p_0_in ),
        .I1(\u1/p_17_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_18_in ),
        .I4(g0_b0_i_71__6_n_0),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_68__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_68__5
       (.I0(key2[33]),
        .I1(roundSel[5]),
        .I2(key3[33]),
        .I3(decrypt),
        .I4(key1[33]),
        .I5(roundSel[4]),
        .O(\u1/p_18_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB4)) 
    g0_b0_i_68__6
       (.I0(roundSel[5]),
        .I1(roundSel[4]),
        .I2(decrypt),
        .O(g0_b0_i_68__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_69
       (.I0(\u1/p_8_in ),
        .I1(\u1/p_9_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_77__5_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_11_in ),
        .O(g0_b0_i_69_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_69__0
       (.I0(g0_b0_i_124_n_0),
        .I1(g0_b0_i_70__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_80__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_85__3_n_0),
        .O(g0_b0_i_69__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_69__1
       (.I0(g0_b0_i_90__3_n_0),
        .I1(g0_b0_i_87__3_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_78__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_102__2_n_0),
        .O(g0_b0_i_69__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_69__2
       (.I0(g0_b0_i_98__0_n_0),
        .I1(roundSel[0]),
        .I2(g0_b0_i_71__4_n_0),
        .I3(decrypt),
        .I4(g0_b0_i_99__0_n_0),
        .O(g0_b0_i_69__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_69__3
       (.I0(\u1/p_3_in ),
        .I1(g0_b0_i_96__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_74__6_n_0),
        .I4(\u1/p_2_in ),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_69__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_69__4
       (.I0(\u1/p_17_in ),
        .I1(\u1/p_18_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_0_in ),
        .I4(g0_b0_i_67__6_n_0),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_69__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_69__5
       (.I0(key2[30]),
        .I1(roundSel[5]),
        .I2(key3[30]),
        .I3(decrypt),
        .I4(key1[30]),
        .I5(roundSel[4]),
        .O(g0_b0_i_69__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_69__6
       (.I0(key2[41]),
        .I1(roundSel[5]),
        .I2(key3[41]),
        .I3(decrypt),
        .I4(key1[41]),
        .I5(roundSel[4]),
        .O(\u1/p_7_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_6__0
       (.I0(desOut[27]),
        .I1(g0_b0_i_22__1_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_23__0_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_24__0_n_0),
        .O(\u0/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_6__1
       (.I0(desOut[59]),
        .I1(g0_b0_i_22__0_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_23__1_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_24__1_n_0),
        .O(\u0/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_6__2
       (.I0(desOut[61]),
        .I1(g0_b0_i_22__2_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_23__2_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_24__2_n_0),
        .O(\u0/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_6__3
       (.I0(desOut[29]),
        .I1(g0_b0_i_22__3_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_23__3_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_24__3_n_0),
        .O(\u0/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_6__4
       (.I0(desOut[63]),
        .I1(g0_b0_i_22__4_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_23__6_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_24__6_n_0),
        .O(\u0/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_6__5
       (.I0(desOut[57]),
        .I1(g0_b0_i_22__6_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_23__4_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_24__4_n_0),
        .O(\u0/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    g0_b0_i_6__6
       (.I0(desOut[31]),
        .I1(g0_b0_i_22__5_n_0),
        .I2(roundSel[3]),
        .I3(g0_b0_i_23__5_n_0),
        .I4(roundSel[2]),
        .I5(g0_b0_i_24__5_n_0),
        .O(\u0/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_7
       (.I0(g0_b0_i_25_n_0),
        .I1(g0_b0_i_26__0_n_0),
        .O(g0_b0_i_7_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_70
       (.I0(\u1/p_1_in ),
        .I1(g0_b0_i_72__5_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_5_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_19_in ),
        .O(g0_b0_i_70_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_70__0
       (.I0(\u1/p_15_in ),
        .I1(g0_b0_i_89__3_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_95__2_n_0),
        .I4(\u1/p_10_in ),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_70__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_70__1
       (.I0(\u1/p_7_in ),
        .I1(g0_b0_i_72__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_71__6_n_0),
        .I4(\u1/p_5_in ),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_70__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_70__2
       (.I0(g0_b0_i_98__2_n_0),
        .I1(g0_b0_i_89__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_100__1_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_86__2_n_0),
        .O(g0_b0_i_70__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_70__3
       (.I0(g0_b0_i_98_n_0),
        .I1(roundSel[0]),
        .I2(g0_b0_i_99_n_0),
        .I3(decrypt),
        .I4(g0_b0_i_72__4_n_0),
        .O(g0_b0_i_70__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_70__4
       (.I0(key1[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_78__6_n_0),
        .I3(roundSel[4]),
        .I4(key3[0]),
        .O(g0_b0_i_70__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_70__5
       (.I0(key2[18]),
        .I1(roundSel[5]),
        .I2(key3[18]),
        .I3(decrypt),
        .I4(key1[18]),
        .I5(roundSel[4]),
        .O(\u1/p_16_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_70__6
       (.I0(key2[36]),
        .I1(roundSel[5]),
        .I2(key3[36]),
        .I3(decrypt),
        .I4(key1[36]),
        .I5(roundSel[4]),
        .O(g0_b0_i_70__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_71
       (.I0(\u1/p_17_in ),
        .I1(\u1/p_3_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_67__6_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_16_in ),
        .O(g0_b0_i_71_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_71__0
       (.I0(g0_b0_i_73__5_n_0),
        .I1(\u1/p_3_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_75__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_16_in ),
        .O(g0_b0_i_71__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_71__1
       (.I0(\u1/p_2_in ),
        .I1(g0_b0_i_98__1_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_96__2_n_0),
        .I4(\u1/p_13_in ),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_71__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_71__2
       (.I0(g0_b0_i_66__5_n_0),
        .I1(g0_b0_i_110__0_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_73__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_67__5_n_0),
        .O(g0_b0_i_71__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_71__3
       (.I0(g0_b0_i_119_n_0),
        .I1(g0_b0_i_66__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_99__1_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_69__5_n_0),
        .O(g0_b0_i_71__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFB08)) 
    g0_b0_i_71__4
       (.I0(key2[0]),
        .I1(roundSel[4]),
        .I2(roundSel[5]),
        .I3(g0_b0_i_78__6_n_0),
        .O(g0_b0_i_71__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_71__5
       (.I0(key2[45]),
        .I1(roundSel[5]),
        .I2(key3[45]),
        .I3(decrypt),
        .I4(key1[45]),
        .I5(roundSel[4]),
        .O(g0_b0_i_71__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_71__6
       (.I0(key2[55]),
        .I1(roundSel[5]),
        .I2(key3[55]),
        .I3(decrypt),
        .I4(key1[55]),
        .I5(roundSel[4]),
        .O(g0_b0_i_71__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_72
       (.I0(g0_b0_i_100__1_n_0),
        .I1(g0_b0_i_80__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_124_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_90__3_n_0),
        .O(g0_b0_i_72_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_72__0
       (.I0(g0_b0_i_124_n_0),
        .I1(\u1/decrypt_int__2 ),
        .I2(g0_b0_i_90__3_n_0),
        .O(g0_b0_i_72__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_72__1
       (.I0(\u1/p_7_in ),
        .I1(\u1/p_14_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_71__6_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(g0_b0_i_74__6_n_0),
        .O(g0_b0_i_72__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_72__2
       (.I0(\u1/p_1_in ),
        .I1(\u1/p_18_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_19_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_0_in ),
        .O(g0_b0_i_72__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_72__3
       (.I0(\u1/p_8_in ),
        .I1(\u1/p_14_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_11_in ),
        .I4(g0_b0_i_74__6_n_0),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_72__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFB08)) 
    g0_b0_i_72__4
       (.I0(key2[0]),
        .I1(roundSel[4]),
        .I2(roundSel[5]),
        .I3(g0_b0_i_72__6_n_0),
        .O(g0_b0_i_72__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_72__5
       (.I0(key2[4]),
        .I1(roundSel[5]),
        .I2(key3[4]),
        .I3(decrypt),
        .I4(key1[4]),
        .I5(roundSel[4]),
        .O(g0_b0_i_72__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_72__6
       (.I0(key2[50]),
        .I1(roundSel[5]),
        .I2(key3[50]),
        .I3(decrypt),
        .I4(key1[50]),
        .I5(roundSel[4]),
        .O(g0_b0_i_72__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_73
       (.I0(g0_b0_i_110__0_n_0),
        .I1(g0_b0_i_73__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_66__5_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_119_n_0),
        .O(g0_b0_i_73_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_73__0
       (.I0(\u1/p_7_in ),
        .I1(g0_b0_i_98__1_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_13_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(g0_b0_i_71__6_n_0),
        .O(g0_b0_i_73__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_73__1
       (.I0(\u1/p_19_in ),
        .I1(\u1/p_16_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_72__5_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_2_in ),
        .O(g0_b0_i_73__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_73__2
       (.I0(g0_b0_i_99__1_n_0),
        .I1(g0_b0_i_115_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_98__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_77__6_n_0),
        .O(g0_b0_i_73__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_73__3
       (.I0(g0_b0_i_73__5_n_0),
        .I1(\u1/p_9_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_75__6_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(g0_b0_i_77__5_n_0),
        .O(g0_b0_i_73__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_73__4
       (.I0(key3[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_72__6_n_0),
        .I3(roundSel[4]),
        .I4(key1[0]),
        .O(g0_b0_i_73__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_73__5
       (.I0(key2[13]),
        .I1(roundSel[5]),
        .I2(key3[13]),
        .I3(decrypt),
        .I4(key1[13]),
        .I5(roundSel[4]),
        .O(g0_b0_i_73__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_73__6
       (.I0(key2[31]),
        .I1(roundSel[5]),
        .I2(key3[31]),
        .I3(decrypt),
        .I4(key1[31]),
        .I5(roundSel[4]),
        .O(g0_b0_i_73__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_74
       (.I0(g0_b0_i_77__5_n_0),
        .I1(g0_b0_i_73__5_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_11_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_9_in ),
        .O(g0_b0_i_74_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    g0_b0_i_74__0
       (.I0(g0_b0_i_79__4_n_0),
        .I1(decrypt),
        .I2(g0_b0_i_100__0_n_0),
        .I3(roundSel[0]),
        .I4(g0_b0_i_101__0_n_0),
        .O(g0_b0_i_74__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_74__1
       (.I0(g0_b0_i_67__6_n_0),
        .I1(g0_b0_i_74__6_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_1_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_3_in ),
        .O(g0_b0_i_74__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_74__2
       (.I0(g0_b0_i_73__5_n_0),
        .I1(\u1/p_18_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_75__6_n_0),
        .I4(\u1/p_0_in ),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_74__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_74__3
       (.I0(g0_b0_i_110__0_n_0),
        .I1(g0_b0_i_102__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_119_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_101__2_n_0),
        .O(g0_b0_i_74__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_74__4
       (.I0(g0_b0_i_65__4_n_0),
        .I1(\u1/decrypt_int__2 ),
        .I2(g0_b0_i_71__5_n_0),
        .O(g0_b0_i_74__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_74__5
       (.I0(g0_b0_i_88__3_n_0),
        .I1(g0_b0_i_68__6_n_0),
        .I2(g0_b0_i_124_n_0),
        .O(g0_b0_i_74__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_74__6
       (.I0(key2[46]),
        .I1(roundSel[5]),
        .I2(key3[46]),
        .I3(decrypt),
        .I4(key1[46]),
        .I5(roundSel[4]),
        .O(g0_b0_i_74__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_75
       (.I0(g0_b0_i_69__5_n_0),
        .I1(g0_b0_i_119_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_110__0_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_66__5_n_0),
        .O(g0_b0_i_75_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_75__0
       (.I0(g0_b0_i_74__6_n_0),
        .I1(\u1/p_7_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_14_in ),
        .I4(g0_b0_i_75__6_n_0),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_75__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_75__1
       (.I0(g0_b0_i_70__6_n_0),
        .I1(g0_b0_i_80__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_72__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_124_n_0),
        .O(g0_b0_i_75__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_75__2
       (.I0(\u1/p_8_in ),
        .I1(g0_b0_i_72__5_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_11_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_5_in ),
        .O(g0_b0_i_75__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_75__3
       (.I0(g0_b0_i_71__6_n_0),
        .I1(g0_b0_i_77__5_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_17_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_14_in ),
        .O(g0_b0_i_75__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_75__4
       (.I0(g0_b0_i_65__4_n_0),
        .I1(g0_b0_i_86__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_67__5_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_87__3_n_0),
        .O(g0_b0_i_75__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFB08)) 
    g0_b0_i_75__5
       (.I0(key2[0]),
        .I1(roundSel[4]),
        .I2(roundSel[5]),
        .I3(g0_b0_i_85__3_n_0),
        .O(g0_b0_i_75__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_75__6
       (.I0(key2[27]),
        .I1(roundSel[5]),
        .I2(key3[27]),
        .I3(decrypt),
        .I4(key1[27]),
        .I5(roundSel[4]),
        .O(g0_b0_i_75__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_76
       (.I0(g0_b0_i_66__5_n_0),
        .I1(g0_b0_i_99__1_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_119_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_73__6_n_0),
        .O(g0_b0_i_76_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_76__0
       (.I0(g0_b0_i_86__2_n_0),
        .I1(g0_b0_i_98__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_89__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_99__1_n_0),
        .O(g0_b0_i_76__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_76__1
       (.I0(\u1/p_16_in ),
        .I1(\u1/p_17_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_3_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(g0_b0_i_71__6_n_0),
        .O(g0_b0_i_76__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_76__2
       (.I0(g0_b0_i_88__3_n_0),
        .I1(g0_b0_i_115_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_85__3_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_77__6_n_0),
        .O(g0_b0_i_76__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_76__3
       (.I0(\u1/p_15_in ),
        .I1(\u1/p_3_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_95__2_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_16_in ),
        .O(g0_b0_i_76__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_76__4
       (.I0(g0_b0_i_75__6_n_0),
        .I1(\u1/p_10_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_7_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_9_in ),
        .O(g0_b0_i_76__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_76__5
       (.I0(key3[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_85__3_n_0),
        .I3(roundSel[4]),
        .I4(key1[0]),
        .O(g0_b0_i_76__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_76__6
       (.I0(key2[32]),
        .I1(roundSel[5]),
        .I2(key3[32]),
        .I3(decrypt),
        .I4(key1[32]),
        .I5(roundSel[4]),
        .O(\u1/p_3_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_77
       (.I0(\u1/p_9_in ),
        .I1(g0_b0_i_75__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_73__5_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_10_in ),
        .O(g0_b0_i_77_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_77__0
       (.I0(g0_b0_i_75__6_n_0),
        .I1(\u1/p_13_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_89__3_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_7_in ),
        .O(g0_b0_i_77__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_77__1
       (.I0(g0_b0_i_89__2_n_0),
        .I1(g0_b0_i_100__1_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_69__5_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_98__2_n_0),
        .O(g0_b0_i_77__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_77__2
       (.I0(g0_b0_i_102__2_n_0),
        .I1(g0_b0_i_90__3_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_87__3_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_100__1_n_0),
        .O(g0_b0_i_77__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_77__3
       (.I0(\u1/p_5_in ),
        .I1(\u1/p_1_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_72__5_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(g0_b0_i_67__6_n_0),
        .O(g0_b0_i_77__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_77__4
       (.I0(g0_b0_i_71__5_n_0),
        .I1(\u1/decrypt_int__2 ),
        .I2(g0_b0_i_67__5_n_0),
        .O(g0_b0_i_77__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_77__5
       (.I0(key2[17]),
        .I1(roundSel[5]),
        .I2(key3[17]),
        .I3(decrypt),
        .I4(key1[17]),
        .I5(roundSel[4]),
        .O(g0_b0_i_77__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_77__6
       (.I0(key2[42]),
        .I1(roundSel[5]),
        .I2(key3[42]),
        .I3(decrypt),
        .I4(key1[42]),
        .I5(roundSel[4]),
        .O(g0_b0_i_77__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_78
       (.I0(g0_b0_i_98__1_n_0),
        .I1(g0_b0_i_67__6_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_17_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_0_in ),
        .O(g0_b0_i_78_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_78__0
       (.I0(\u1/p_14_in ),
        .I1(g0_b0_i_71__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_77__5_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_7_in ),
        .O(g0_b0_i_78__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_78__1
       (.I0(\u1/p_11_in ),
        .I1(\u1/p_0_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_73__5_n_0),
        .I4(g0_b0_i_98__1_n_0),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_78__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_78__2
       (.I0(g0_b0_i_87__3_n_0),
        .I1(g0_b0_i_78__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_86__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_90__3_n_0),
        .O(g0_b0_i_78__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_78__3
       (.I0(g0_b0_i_115_n_0),
        .I1(g0_b0_i_79__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_101__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_78__6_n_0),
        .O(g0_b0_i_78__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_78__4
       (.I0(key1[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_65__4_n_0),
        .I3(roundSel[4]),
        .I4(key3[0]),
        .O(g0_b0_i_78__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_78__5
       (.I0(key2[10]),
        .I1(roundSel[5]),
        .I2(key3[10]),
        .I3(decrypt),
        .I4(key1[10]),
        .I5(roundSel[4]),
        .O(\u1/p_8_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_78__6
       (.I0(key2[35]),
        .I1(roundSel[5]),
        .I2(key3[35]),
        .I3(decrypt),
        .I4(key1[35]),
        .I5(roundSel[4]),
        .O(g0_b0_i_78__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_79
       (.I0(g0_b0_i_102__2_n_0),
        .I1(g0_b0_i_72__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_70__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_87__3_n_0),
        .O(g0_b0_i_79_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_79__0
       (.I0(g0_b0_i_89__3_n_0),
        .I1(\u1/p_19_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_13_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_1_in ),
        .O(g0_b0_i_79__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_79__1
       (.I0(\u1/p_3_in ),
        .I1(g0_b0_i_67__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_74__6_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_17_in ),
        .O(g0_b0_i_79__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_79__2
       (.I0(g0_b0_i_95__2_n_0),
        .I1(\u1/p_5_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_8_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_18_in ),
        .O(g0_b0_i_79__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_79__3
       (.I0(g0_b0_i_101__2_n_0),
        .I1(g0_b0_i_88__3_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_102__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_79__6_n_0),
        .O(g0_b0_i_79__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFB08)) 
    g0_b0_i_79__4
       (.I0(key2[0]),
        .I1(roundSel[4]),
        .I2(roundSel[5]),
        .I3(g0_b0_i_65__4_n_0),
        .O(g0_b0_i_79__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_79__5
       (.I0(key2[24]),
        .I1(roundSel[5]),
        .I2(key3[24]),
        .I3(decrypt),
        .I4(key1[24]),
        .I5(roundSel[4]),
        .O(\u1/p_11_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_79__6
       (.I0(key2[49]),
        .I1(roundSel[5]),
        .I2(key3[49]),
        .I3(decrypt),
        .I4(key1[49]),
        .I5(roundSel[4]),
        .O(g0_b0_i_79__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_7__0
       (.I0(g0_b0_i_25__0_n_0),
        .I1(g0_b0_i_26__1_n_0),
        .O(g0_b0_i_7__0_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_7__1
       (.I0(g0_b0_i_25__1_n_0),
        .I1(g0_b0_i_26__2_n_0),
        .O(g0_b0_i_7__1_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_7__2
       (.I0(g0_b0_i_25__2_n_0),
        .I1(g0_b0_i_26__3_n_0),
        .O(g0_b0_i_7__2_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_7__3
       (.I0(g0_b0_i_25__3_n_0),
        .I1(g0_b0_i_26__4_n_0),
        .O(g0_b0_i_7__3_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_7__4
       (.I0(g0_b0_i_25__4_n_0),
        .I1(g0_b0_i_26__5_n_0),
        .O(g0_b0_i_7__4_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_7__5
       (.I0(g0_b0_i_25__5_n_0),
        .I1(g0_b0_i_26__6_n_0),
        .O(g0_b0_i_7__5_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 g0_b0_i_7__6
       (.I0(g0_b0_i_25__6_n_0),
        .I1(g0_b0_i_26_n_0),
        .O(g0_b0_i_7__6_n_0),
        .S(roundSel[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_8
       (.I0(g0_b0_i_27_n_0),
        .I1(g0_b0_i_28__0_n_0),
        .O(g0_b0_i_8_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_80
       (.I0(g0_b0_i_101__2_n_0),
        .I1(g0_b0_i_70__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_85__3_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_102__2_n_0),
        .O(g0_b0_i_80_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    g0_b0_i_80__0
       (.I0(g0_b0_i_86__1_n_0),
        .I1(decrypt),
        .I2(g0_b0_i_93__3_n_0),
        .I3(roundSel[0]),
        .I4(g0_b0_i_94__0_n_0),
        .O(g0_b0_i_80__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_80__1
       (.I0(g0_b0_i_115_n_0),
        .I1(g0_b0_i_67__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_101__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_65__4_n_0),
        .O(g0_b0_i_80__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_80__2
       (.I0(\u1/p_9_in ),
        .I1(g0_b0_i_96__2_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_10_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_2_in ),
        .O(g0_b0_i_80__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_80__3
       (.I0(g0_b0_i_72__5_n_0),
        .I1(\u1/p_19_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_16_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_1_in ),
        .O(g0_b0_i_80__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_80__4
       (.I0(g0_b0_i_96__2_n_0),
        .I1(\u1/p_16_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_15_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_72__5_n_0),
        .O(g0_b0_i_80__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_80__5
       (.I0(key2[3]),
        .I1(roundSel[5]),
        .I2(key3[3]),
        .I3(decrypt),
        .I4(key1[3]),
        .I5(roundSel[4]),
        .O(\u1/p_14_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_80__6
       (.I0(key2[28]),
        .I1(roundSel[5]),
        .I2(key3[28]),
        .I3(decrypt),
        .I4(key1[28]),
        .I5(roundSel[4]),
        .O(g0_b0_i_80__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_81
       (.I0(\u1/p_5_in ),
        .I1(\u1/p_2_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_19_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(g0_b0_i_72__5_n_0),
        .O(g0_b0_i_81_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_81__0
       (.I0(\u1/p_10_in ),
        .I1(\u1/p_7_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_75__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_89__3_n_0),
        .O(g0_b0_i_81__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_81__1
       (.I0(\u1/p_18_in ),
        .I1(\u1/p_19_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_1_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_5_in ),
        .O(g0_b0_i_81__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_81__2
       (.I0(g0_b0_i_127_n_0),
        .I1(roundSel[0]),
        .I2(g0_b0_i_92__3_n_0),
        .I3(decrypt),
        .I4(g0_b0_i_84__6_n_0),
        .O(g0_b0_i_81__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_81__3
       (.I0(g0_b0_i_77__6_n_0),
        .I1(g0_b0_i_65__4_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_115_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_72__6_n_0),
        .O(g0_b0_i_81__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_81__4
       (.I0(g0_b0_i_110__0_n_0),
        .I1(g0_b0_i_80__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_119_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_124_n_0),
        .O(g0_b0_i_81__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_81__5
       (.I0(g0_b0_i_80__6_n_0),
        .I1(g0_b0_i_119_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_77__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_110__0_n_0),
        .O(g0_b0_i_81__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_81__6
       (.I0(\u1/p_14_in ),
        .I1(g0_b0_i_95__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_77__5_n_0),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_15_in ),
        .O(g0_b0_i_81__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_82
       (.I0(g0_b0_i_73__5_n_0),
        .I1(g0_b0_i_89__3_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_10_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(g0_b0_i_75__6_n_0),
        .O(g0_b0_i_82_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_82__0
       (.I0(g0_b0_i_66__5_n_0),
        .I1(g0_b0_i_78__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_73__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_90__3_n_0),
        .O(g0_b0_i_82__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_82__1
       (.I0(\u1/p_0_in ),
        .I1(\u1/p_15_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_18_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(g0_b0_i_96__2_n_0),
        .O(g0_b0_i_82__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_82__2
       (.I0(g0_b0_i_77__5_n_0),
        .I1(\u1/p_17_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_9_in ),
        .I4(g0_b0_i_71__6_n_0),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_82__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_82__3
       (.I0(g0_b0_i_124_n_0),
        .I1(g0_b0_i_110__0_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_80__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_67__5_n_0),
        .O(g0_b0_i_82__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_82__4
       (.I0(g0_b0_i_65__4_n_0),
        .I1(g0_b0_i_115_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_67__5_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_77__6_n_0),
        .O(g0_b0_i_82__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    g0_b0_i_82__5
       (.I0(g0_b0_i_91__3_n_0),
        .I1(decrypt),
        .I2(g0_b0_i_92__3_n_0),
        .I3(roundSel[0]),
        .I4(g0_b0_i_100_n_0),
        .O(g0_b0_i_82__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_82__6
       (.I0(g0_b0_i_98__1_n_0),
        .I1(g0_b0_i_96__2_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_0_in ),
        .I4(\u1/p_2_in ),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_82__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_83
       (.I0(\u1/p_8_in ),
        .I1(g0_b0_i_98__1_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_11_in ),
        .I4(g0_b0_i_65__6_n_0),
        .I5(\u1/p_13_in ),
        .O(g0_b0_i_83_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_83__0
       (.I0(g0_b0_i_89__2_n_0),
        .I1(g0_b0_i_88__3_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_69__5_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_79__6_n_0),
        .O(g0_b0_i_83__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_83__1
       (.I0(g0_b0_i_74__6_n_0),
        .I1(\u1/p_1_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_14_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_67__6_n_0),
        .O(g0_b0_i_83__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_83__2
       (.I0(\u1/p_13_in ),
        .I1(\u1/p_8_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_98__1_n_0),
        .I4(g0_b0_i_95__2_n_0),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_83__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_83__3
       (.I0(g0_b0_i_70__6_n_0),
        .I1(g0_b0_i_102__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_72__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_101__2_n_0),
        .O(g0_b0_i_83__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_83__4
       (.I0(g0_b0_i_102__0_n_0),
        .I1(roundSel[0]),
        .I2(g0_b0_i_103__1_n_0),
        .I3(decrypt),
        .I4(g0_b0_i_84__5_n_0),
        .O(g0_b0_i_83__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_83__5
       (.I0(g0_b0_i_99__1_n_0),
        .I1(\u1/decrypt_int__2 ),
        .I2(g0_b0_i_124_n_0),
        .O(g0_b0_i_83__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_83__6
       (.I0(g0_b0_i_89__3_n_0),
        .I1(g0_b0_i_95__2_n_0),
        .I2(roundSel[0]),
        .I3(\u1/p_13_in ),
        .I4(\u1/p_15_in ),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_83__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_84
       (.I0(\u1/p_15_in ),
        .I1(\u1/p_18_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_95__2_n_0),
        .I4(\u1/p_0_in ),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_84_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_84__0
       (.I0(g0_b0_i_87__3_n_0),
        .I1(g0_b0_i_70__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_86__2_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_85__3_n_0),
        .O(g0_b0_i_84__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_84__1
       (.I0(\u1/p_16_in ),
        .I1(\u1/p_2_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_3_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_19_in ),
        .O(g0_b0_i_84__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_84__2
       (.I0(g0_b0_i_98__2_n_0),
        .I1(\u1/decrypt_int__2 ),
        .I2(g0_b0_i_71__5_n_0),
        .O(g0_b0_i_84__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_84__3
       (.I0(\u1/p_10_in ),
        .I1(g0_b0_i_73__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_89__3_n_0),
        .I4(\u1/p_11_in ),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_84__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_84__4
       (.I0(\u1/p_9_in ),
        .I1(\u1/p_11_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_10_in ),
        .I4(\u1/p_8_in ),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_84__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFB08)) 
    g0_b0_i_84__5
       (.I0(key2[0]),
        .I1(roundSel[4]),
        .I2(roundSel[5]),
        .I3(g0_b0_i_119_n_0),
        .O(g0_b0_i_84__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_84__6
       (.I0(key3[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_98__2_n_0),
        .I3(roundSel[4]),
        .I4(key1[0]),
        .O(g0_b0_i_84__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_85
       (.I0(g0_b0_i_124_n_0),
        .I1(g0_b0_i_78__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_90__3_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_80__6_n_0),
        .O(g0_b0_i_85_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_85__0
       (.I0(\u1/p_2_in ),
        .I1(g0_b0_i_72__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_96__2_n_0),
        .I4(\u1/p_5_in ),
        .I5(g0_b0_i_65__6_n_0),
        .O(g0_b0_i_85__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_85__1
       (.I0(key3[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_119_n_0),
        .I3(roundSel[4]),
        .I4(key1[0]),
        .O(g0_b0_i_85__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_85__2
       (.I0(key1[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_99__1_n_0),
        .I3(roundSel[4]),
        .I4(key3[0]),
        .O(g0_b0_i_85__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_85__3
       (.I0(key2[22]),
        .I1(roundSel[5]),
        .I2(key3[22]),
        .I3(decrypt),
        .I4(key1[22]),
        .I5(roundSel[4]),
        .O(g0_b0_i_85__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_85__4
       (.I0(key2[54]),
        .I1(roundSel[5]),
        .I2(key3[54]),
        .I3(decrypt),
        .I4(key1[54]),
        .I5(roundSel[4]),
        .O(\u1/p_19_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_86
       (.I0(g0_b0_i_101__1_n_0),
        .I1(roundSel[0]),
        .I2(g0_b0_i_102__1_n_0),
        .I3(decrypt),
        .I4(g0_b0_i_89__1_n_0),
        .O(g0_b0_i_86_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_86__0
       (.I0(g0_b0_i_99__1_n_0),
        .I1(\u1/decrypt_int__2 ),
        .I2(g0_b0_i_71__5_n_0),
        .O(g0_b0_i_86__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFB08)) 
    g0_b0_i_86__1
       (.I0(key2[0]),
        .I1(roundSel[4]),
        .I2(roundSel[5]),
        .I3(g0_b0_i_99__1_n_0),
        .O(g0_b0_i_86__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_86__2
       (.I0(key2[2]),
        .I1(roundSel[5]),
        .I2(key3[2]),
        .I3(decrypt),
        .I4(key1[2]),
        .I5(roundSel[4]),
        .O(g0_b0_i_86__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_86__3
       (.I0(key2[11]),
        .I1(roundSel[5]),
        .I2(key3[11]),
        .I3(decrypt),
        .I4(key1[11]),
        .I5(roundSel[4]),
        .O(\u1/p_2_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_87
       (.I0(g0_b0_i_89__2_n_0),
        .I1(g0_b0_i_110__0_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_67__5_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_69__5_n_0),
        .O(g0_b0_i_87_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_87__0
       (.I0(g0_b0_i_85__3_n_0),
        .I1(g0_b0_i_87__3_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_102__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_70__6_n_0),
        .O(g0_b0_i_87__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_87__1
       (.I0(g0_b0_i_66__5_n_0),
        .I1(g0_b0_i_70__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_73__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_85__3_n_0),
        .O(g0_b0_i_87__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_87__2
       (.I0(key2[40]),
        .I1(roundSel[5]),
        .I2(key3[40]),
        .I3(decrypt),
        .I4(key1[40]),
        .I5(roundSel[4]),
        .O(\u1/p_1_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_87__3
       (.I0(key2[43]),
        .I1(roundSel[5]),
        .I2(key3[43]),
        .I3(decrypt),
        .I4(key1[43]),
        .I5(roundSel[4]),
        .O(g0_b0_i_87__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_88
       (.I0(g0_b0_i_87__3_n_0),
        .I1(g0_b0_i_99__1_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_86__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_119_n_0),
        .O(g0_b0_i_88_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_88__0
       (.I0(g0_b0_i_79__6_n_0),
        .I1(g0_b0_i_89__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_88__3_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_86__2_n_0),
        .O(g0_b0_i_88__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_88__1
       (.I0(g0_b0_i_89__2_n_0),
        .I1(g0_b0_i_65__4_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_69__5_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_72__6_n_0),
        .O(g0_b0_i_88__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_88__2
       (.I0(key2[6]),
        .I1(roundSel[5]),
        .I2(key3[6]),
        .I3(decrypt),
        .I4(key1[6]),
        .I5(roundSel[4]),
        .O(\u1/p_9_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_88__3
       (.I0(key2[8]),
        .I1(roundSel[5]),
        .I2(key3[8]),
        .I3(decrypt),
        .I4(key1[8]),
        .I5(roundSel[4]),
        .O(g0_b0_i_88__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_89
       (.I0(g0_b0_i_101__2_n_0),
        .I1(g0_b0_i_100__1_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_102__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_98__2_n_0),
        .O(g0_b0_i_89_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_89__0
       (.I0(g0_b0_i_90__3_n_0),
        .I1(g0_b0_i_66__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_78__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_69__5_n_0),
        .O(g0_b0_i_89__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFB08)) 
    g0_b0_i_89__1
       (.I0(key2[0]),
        .I1(roundSel[4]),
        .I2(roundSel[5]),
        .I3(g0_b0_i_79__6_n_0),
        .O(g0_b0_i_89__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_89__2
       (.I0(key2[16]),
        .I1(roundSel[5]),
        .I2(key3[16]),
        .I3(decrypt),
        .I4(key1[16]),
        .I5(roundSel[4]),
        .O(g0_b0_i_89__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_89__3
       (.I0(key2[34]),
        .I1(roundSel[5]),
        .I2(key3[34]),
        .I3(decrypt),
        .I4(key1[34]),
        .I5(roundSel[4]),
        .O(g0_b0_i_89__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_8__0
       (.I0(g0_b0_i_27__0_n_0),
        .I1(g0_b0_i_28__5_n_0),
        .O(g0_b0_i_8__0_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_8__1
       (.I0(g0_b0_i_27__1_n_0),
        .I1(g0_b0_i_28__1_n_0),
        .O(g0_b0_i_8__1_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_8__2
       (.I0(g0_b0_i_27__2_n_0),
        .I1(g0_b0_i_28__6_n_0),
        .O(g0_b0_i_8__2_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_8__3
       (.I0(g0_b0_i_27__3_n_0),
        .I1(g0_b0_i_28__3_n_0),
        .O(g0_b0_i_8__3_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_8__4
       (.I0(g0_b0_i_27__4_n_0),
        .I1(g0_b0_i_28__2_n_0),
        .O(g0_b0_i_8__4_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_8__5
       (.I0(g0_b0_i_27__5_n_0),
        .I1(g0_b0_i_28__4_n_0),
        .O(g0_b0_i_8__5_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_8__6
       (.I0(g0_b0_i_27__6_n_0),
        .I1(g0_b0_i_28_n_0),
        .O(g0_b0_i_8__6_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_9
       (.I0(g0_b0_i_29__6_n_0),
        .I1(g0_b0_i_30_n_0),
        .O(g0_b0_i_9_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_90
       (.I0(g0_b0_i_77__6_n_0),
        .I1(g0_b0_i_78__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_115_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_90__3_n_0),
        .O(g0_b0_i_90_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_90__0
       (.I0(g0_b0_i_98__2_n_0),
        .I1(g0_b0_i_71__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_100__1_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_73__6_n_0),
        .O(g0_b0_i_90__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_90__1
       (.I0(key3[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_79__6_n_0),
        .I3(roundSel[4]),
        .I4(key1[0]),
        .O(g0_b0_i_90__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_90__2
       (.I0(key2[20]),
        .I1(roundSel[5]),
        .I2(key3[20]),
        .I3(decrypt),
        .I4(key1[20]),
        .I5(roundSel[4]),
        .O(\u1/p_10_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_90__3
       (.I0(key2[21]),
        .I1(roundSel[5]),
        .I2(key3[21]),
        .I3(decrypt),
        .I4(key1[21]),
        .I5(roundSel[4]),
        .O(g0_b0_i_90__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    g0_b0_i_91
       (.I0(g0_b0_i_104__1_n_0),
        .I1(decrypt),
        .I2(g0_b0_i_96__1_n_0),
        .I3(roundSel[0]),
        .I4(g0_b0_i_105_n_0),
        .O(g0_b0_i_91_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_91__0
       (.I0(\u1/p_0_in ),
        .I1(\u1/p_1_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_67__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(\u1/p_18_in ),
        .O(g0_b0_i_91__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_91__1
       (.I0(g0_b0_i_88__3_n_0),
        .I1(\u1/decrypt_int__2 ),
        .I2(g0_b0_i_71__5_n_0),
        .O(g0_b0_i_91__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_91__2
       (.I0(key3[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_88__3_n_0),
        .I3(roundSel[4]),
        .I4(key1[0]),
        .O(g0_b0_i_91__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_91__3
       (.I0(key1[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_98__2_n_0),
        .I3(roundSel[4]),
        .I4(key3[0]),
        .O(g0_b0_i_91__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_92
       (.I0(g0_b0_i_86__2_n_0),
        .I1(g0_b0_i_67__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_65__4_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_89__2_n_0),
        .O(g0_b0_i_92_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_92__0
       (.I0(g0_b0_i_73__6_n_0),
        .I1(g0_b0_i_79__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_71__5_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_78__6_n_0),
        .O(g0_b0_i_92__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_92__1
       (.I0(\u1/p_13_in ),
        .I1(\u1/p_2_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_98__1_n_0),
        .I4(\u1/p_19_in ),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_92__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_92__2
       (.I0(g0_b0_i_85__3_n_0),
        .I1(\u1/decrypt_int__2 ),
        .I2(g0_b0_i_71__5_n_0),
        .O(g0_b0_i_92__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFB08)) 
    g0_b0_i_92__3
       (.I0(key2[0]),
        .I1(roundSel[4]),
        .I2(roundSel[5]),
        .I3(g0_b0_i_98__2_n_0),
        .O(g0_b0_i_92__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_93
       (.I0(g0_b0_i_102__2_n_0),
        .I1(g0_b0_i_119_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_87__3_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_110__0_n_0),
        .O(g0_b0_i_93_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_93__0
       (.I0(g0_b0_i_69__5_n_0),
        .I1(g0_b0_i_85__3_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_66__5_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_88__3_n_0),
        .O(g0_b0_i_93__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    g0_b0_i_93__1
       (.I0(\u1/p_10_in ),
        .I1(\u1/p_15_in ),
        .I2(roundSel[0]),
        .I3(g0_b0_i_89__3_n_0),
        .I4(g0_b0_i_96__2_n_0),
        .I5(g0_b0_i_68__6_n_0),
        .O(g0_b0_i_93__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_93__2
       (.I0(g0_b0_i_100__1_n_0),
        .I1(g0_b0_i_68__6_n_0),
        .I2(g0_b0_i_71__5_n_0),
        .O(g0_b0_i_93__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_93__3
       (.I0(key3[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_99__1_n_0),
        .I3(roundSel[4]),
        .I4(key1[0]),
        .O(g0_b0_i_93__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_94
       (.I0(g0_b0_i_88__3_n_0),
        .I1(g0_b0_i_102__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_101__2_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_85__3_n_0),
        .O(g0_b0_i_94_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_94__0
       (.I0(g0_b0_i_71__5_n_0),
        .I1(\u1/decrypt_int__2 ),
        .I2(g0_b0_i_98__2_n_0),
        .O(g0_b0_i_94__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_94__1
       (.I0(g0_b0_i_115_n_0),
        .I1(g0_b0_i_98__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_101__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_99__1_n_0),
        .O(g0_b0_i_94__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_94__2
       (.I0(g0_b0_i_86__2_n_0),
        .I1(g0_b0_i_72__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_89__2_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_70__6_n_0),
        .O(g0_b0_i_94__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_94__3
       (.I0(g0_b0_i_77__5_n_0),
        .I1(\u1/p_8_in ),
        .I2(roundSel[0]),
        .I3(\u1/p_9_in ),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_95__2_n_0),
        .O(g0_b0_i_94__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_95
       (.I0(g0_b0_i_78__6_n_0),
        .I1(g0_b0_i_86__2_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_79__6_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_87__3_n_0),
        .O(g0_b0_i_95_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_95__0
       (.I0(g0_b0_i_80__6_n_0),
        .I1(g0_b0_i_90__3_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_77__6_n_0),
        .I4(\u1/decrypt_int__2 ),
        .I5(g0_b0_i_100__1_n_0),
        .O(g0_b0_i_95__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_95__1
       (.I0(g0_b0_i_124_n_0),
        .I1(\u1/decrypt_int__2 ),
        .I2(g0_b0_i_100__1_n_0),
        .O(g0_b0_i_95__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_95__2
       (.I0(key2[53]),
        .I1(roundSel[5]),
        .I2(key3[53]),
        .I3(decrypt),
        .I4(key1[53]),
        .I5(roundSel[4]),
        .O(g0_b0_i_95__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_96
       (.I0(g0_b0_i_98__2_n_0),
        .I1(\u1/decrypt_int__2 ),
        .I2(g0_b0_i_124_n_0),
        .O(g0_b0_i_96_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_96__0
       (.I0(g0_b0_i_100__1_n_0),
        .I1(g0_b0_i_69__5_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_90__3_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_89__2_n_0),
        .O(g0_b0_i_96__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFB08)) 
    g0_b0_i_96__1
       (.I0(key2[0]),
        .I1(roundSel[4]),
        .I2(roundSel[5]),
        .I3(g0_b0_i_90__3_n_0),
        .O(g0_b0_i_96__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_96__2
       (.I0(key2[25]),
        .I1(roundSel[5]),
        .I2(key3[25]),
        .I3(decrypt),
        .I4(key1[25]),
        .I5(roundSel[4]),
        .O(g0_b0_i_96__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    g0_b0_i_97
       (.I0(g0_b0_i_99__1_n_0),
        .I1(g0_b0_i_73__6_n_0),
        .I2(roundSel[0]),
        .I3(g0_b0_i_98__2_n_0),
        .I4(g0_b0_i_68__6_n_0),
        .I5(g0_b0_i_66__5_n_0),
        .O(g0_b0_i_97_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_97__0
       (.I0(key1[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_100__1_n_0),
        .I3(roundSel[4]),
        .I4(key3[0]),
        .O(g0_b0_i_97__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_97__1
       (.I0(key3[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_90__3_n_0),
        .I3(roundSel[4]),
        .I4(key1[0]),
        .O(g0_b0_i_97__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_97__2
       (.I0(key2[39]),
        .I1(roundSel[5]),
        .I2(key3[39]),
        .I3(decrypt),
        .I4(key1[39]),
        .I5(roundSel[4]),
        .O(\u1/p_15_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_98
       (.I0(g0_b0_i_71__5_n_0),
        .I1(\u1/decrypt_int__2 ),
        .I2(g0_b0_i_65__4_n_0),
        .O(g0_b0_i_98_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    g0_b0_i_98__0
       (.I0(g0_b0_i_90__3_n_0),
        .I1(\u1/decrypt_int__2 ),
        .I2(g0_b0_i_124_n_0),
        .O(g0_b0_i_98__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_98__1
       (.I0(key2[5]),
        .I1(roundSel[5]),
        .I2(key3[5]),
        .I3(decrypt),
        .I4(key1[5]),
        .I5(roundSel[4]),
        .O(g0_b0_i_98__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_98__2
       (.I0(key2[52]),
        .I1(roundSel[5]),
        .I2(key3[52]),
        .I3(decrypt),
        .I4(key1[52]),
        .I5(roundSel[4]),
        .O(g0_b0_i_98__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_99
       (.I0(key1[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_72__6_n_0),
        .I3(roundSel[4]),
        .I4(key3[0]),
        .O(g0_b0_i_99_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    g0_b0_i_99__0
       (.I0(key3[0]),
        .I1(roundSel[5]),
        .I2(g0_b0_i_78__6_n_0),
        .I3(roundSel[4]),
        .I4(key1[0]),
        .O(g0_b0_i_99__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_99__1
       (.I0(key2[38]),
        .I1(roundSel[5]),
        .I2(key3[38]),
        .I3(decrypt),
        .I4(key1[38]),
        .I5(roundSel[4]),
        .O(g0_b0_i_99__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAFCF330C0)) 
    g0_b0_i_99__2
       (.I0(key2[48]),
        .I1(roundSel[5]),
        .I2(key3[48]),
        .I3(decrypt),
        .I4(key1[48]),
        .I5(roundSel[4]),
        .O(\u1/p_13_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_9__0
       (.I0(g0_b0_i_29__1_n_0),
        .I1(g0_b0_i_30__0_n_0),
        .O(g0_b0_i_9__0_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_9__1
       (.I0(g0_b0_i_29__0_n_0),
        .I1(g0_b0_i_30__1_n_0),
        .O(g0_b0_i_9__1_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_9__2
       (.I0(g0_b0_i_29__2_n_0),
        .I1(g0_b0_i_30__2_n_0),
        .O(g0_b0_i_9__2_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_9__3
       (.I0(g0_b0_i_29__4_n_0),
        .I1(g0_b0_i_30__3_n_0),
        .O(g0_b0_i_9__3_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_9__4
       (.I0(g0_b0_i_29__3_n_0),
        .I1(g0_b0_i_30__4_n_0),
        .O(g0_b0_i_9__4_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_9__5
       (.I0(g0_b0_i_29__5_n_0),
        .I1(g0_b0_i_30__5_n_0),
        .O(g0_b0_i_9__5_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 g0_b0_i_9__6
       (.I0(g0_b0_i_29_n_0),
        .I1(g0_b0_i_30__6_n_0),
        .O(g0_b0_i_9__6_n_0),
        .S(roundSel[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1
       (.I0(\u0/X [41]),
        .I1(\u0/X [40]),
        .I2(\u0/X [39]),
        .I3(\u0/X [38]),
        .I4(\u0/X [42]),
        .I5(\u0/X [37]),
        .O(out[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__0
       (.I0(\u0/X [17]),
        .I1(\u0/X [16]),
        .I2(\u0/X [15]),
        .I3(\u0/X [14]),
        .I4(\u0/X [18]),
        .I5(\u0/X [13]),
        .O(out[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__1
       (.I0(\u0/X [35]),
        .I1(\u0/X [34]),
        .I2(\u0/X [33]),
        .I3(\u0/X [32]),
        .I4(\u0/X [36]),
        .I5(\u0/X [31]),
        .O(out[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__2
       (.I0(\u0/X [11]),
        .I1(\u0/X [10]),
        .I2(\u0/X [9]),
        .I3(\u0/X [8]),
        .I4(\u0/X [12]),
        .I5(\u0/X [7]),
        .O(out[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__3
       (.I0(\u0/X [47]),
        .I1(\u0/X [46]),
        .I2(\u0/X [45]),
        .I3(\u0/X [44]),
        .I4(\u0/X [48]),
        .I5(\u0/X [43]),
        .O(out[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__4
       (.I0(\u0/X [23]),
        .I1(\u0/X [22]),
        .I2(\u0/X [21]),
        .I3(\u0/X [20]),
        .I4(\u0/X [24]),
        .I5(\u0/X [19]),
        .O(out[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__5
       (.I0(\u0/X [29]),
        .I1(\u0/X [28]),
        .I2(\u0/X [27]),
        .I3(\u0/X [26]),
        .I4(\u0/X [30]),
        .I5(\u0/X [25]),
        .O(out[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__6
       (.I0(\u0/X [5]),
        .I1(\u0/X [4]),
        .I2(\u0/X [3]),
        .I3(\u0/X [2]),
        .I4(\u0/X [6]),
        .I5(\u0/X [1]),
        .O(out[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2
       (.I0(\u0/X [41]),
        .I1(\u0/X [40]),
        .I2(\u0/X [39]),
        .I3(\u0/X [38]),
        .I4(\u0/X [42]),
        .I5(\u0/X [37]),
        .O(out[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__0
       (.I0(\u0/X [17]),
        .I1(\u0/X [16]),
        .I2(\u0/X [15]),
        .I3(\u0/X [14]),
        .I4(\u0/X [18]),
        .I5(\u0/X [13]),
        .O(out[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__1
       (.I0(\u0/X [35]),
        .I1(\u0/X [34]),
        .I2(\u0/X [33]),
        .I3(\u0/X [32]),
        .I4(\u0/X [36]),
        .I5(\u0/X [31]),
        .O(out[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__2
       (.I0(\u0/X [11]),
        .I1(\u0/X [10]),
        .I2(\u0/X [9]),
        .I3(\u0/X [8]),
        .I4(\u0/X [12]),
        .I5(\u0/X [7]),
        .O(out[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__3
       (.I0(\u0/X [47]),
        .I1(\u0/X [46]),
        .I2(\u0/X [45]),
        .I3(\u0/X [44]),
        .I4(\u0/X [48]),
        .I5(\u0/X [43]),
        .O(out[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__4
       (.I0(\u0/X [23]),
        .I1(\u0/X [22]),
        .I2(\u0/X [21]),
        .I3(\u0/X [20]),
        .I4(\u0/X [24]),
        .I5(\u0/X [19]),
        .O(out[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__5
       (.I0(\u0/X [29]),
        .I1(\u0/X [28]),
        .I2(\u0/X [27]),
        .I3(\u0/X [26]),
        .I4(\u0/X [30]),
        .I5(\u0/X [25]),
        .O(out[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__6
       (.I0(\u0/X [5]),
        .I1(\u0/X [4]),
        .I2(\u0/X [3]),
        .I3(\u0/X [2]),
        .I4(\u0/X [6]),
        .I5(\u0/X [1]),
        .O(out[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3
       (.I0(\u0/X [41]),
        .I1(\u0/X [40]),
        .I2(\u0/X [39]),
        .I3(\u0/X [38]),
        .I4(\u0/X [42]),
        .I5(\u0/X [37]),
        .O(out[32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__0
       (.I0(\u0/X [17]),
        .I1(\u0/X [16]),
        .I2(\u0/X [15]),
        .I3(\u0/X [14]),
        .I4(\u0/X [18]),
        .I5(\u0/X [13]),
        .O(out[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__1
       (.I0(\u0/X [35]),
        .I1(\u0/X [34]),
        .I2(\u0/X [33]),
        .I3(\u0/X [32]),
        .I4(\u0/X [36]),
        .I5(\u0/X [31]),
        .O(out[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__2
       (.I0(\u0/X [11]),
        .I1(\u0/X [10]),
        .I2(\u0/X [9]),
        .I3(\u0/X [8]),
        .I4(\u0/X [12]),
        .I5(\u0/X [7]),
        .O(out[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__3
       (.I0(\u0/X [47]),
        .I1(\u0/X [46]),
        .I2(\u0/X [45]),
        .I3(\u0/X [44]),
        .I4(\u0/X [48]),
        .I5(\u0/X [43]),
        .O(out[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__4
       (.I0(\u0/X [23]),
        .I1(\u0/X [22]),
        .I2(\u0/X [21]),
        .I3(\u0/X [20]),
        .I4(\u0/X [24]),
        .I5(\u0/X [19]),
        .O(out[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__5
       (.I0(\u0/X [29]),
        .I1(\u0/X [28]),
        .I2(\u0/X [27]),
        .I3(\u0/X [26]),
        .I4(\u0/X [30]),
        .I5(\u0/X [25]),
        .O(out[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__6
       (.I0(\u0/X [5]),
        .I1(\u0/X [4]),
        .I2(\u0/X [3]),
        .I3(\u0/X [2]),
        .I4(\u0/X [6]),
        .I5(\u0/X [1]),
        .O(out[9]));
endmodule
