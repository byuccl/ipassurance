module ahbctrl
   (rst,
    clk,
    \msti[hgrant] ,
    \msti[hready] ,
    \msti[hresp] ,
    \msti[hrdata] ,
    \msti[hirq] ,
    \msti[testen] ,
    \msti[testrst] ,
    \msti[scanen] ,
    \msti[testoen] ,
    \msti[testin] ,
    \msto[15][hbusreq] ,
    \msto[15][hlock] ,
    \msto[15][htrans] ,
    \msto[15][haddr] ,
    \msto[15][hwrite] ,
    \msto[15][hsize] ,
    \msto[15][hburst] ,
    \msto[15][hprot] ,
    \msto[15][hwdata] ,
    \msto[15][hirq] ,
    \msto[15][hconfig][0] ,
    \msto[15][hconfig][1] ,
    \msto[15][hconfig][2] ,
    \msto[15][hconfig][3] ,
    \msto[15][hconfig][4] ,
    \msto[15][hconfig][5] ,
    \msto[15][hconfig][6] ,
    \msto[15][hconfig][7] ,
    \msto[15][hindex] ,
    \msto[14][hbusreq] ,
    \msto[14][hlock] ,
    \msto[14][htrans] ,
    \msto[14][haddr] ,
    \msto[14][hwrite] ,
    \msto[14][hsize] ,
    \msto[14][hburst] ,
    \msto[14][hprot] ,
    \msto[14][hwdata] ,
    \msto[14][hirq] ,
    \msto[14][hconfig][0] ,
    \msto[14][hconfig][1] ,
    \msto[14][hconfig][2] ,
    \msto[14][hconfig][3] ,
    \msto[14][hconfig][4] ,
    \msto[14][hconfig][5] ,
    \msto[14][hconfig][6] ,
    \msto[14][hconfig][7] ,
    \msto[14][hindex] ,
    \msto[13][hbusreq] ,
    \msto[13][hlock] ,
    \msto[13][htrans] ,
    \msto[13][haddr] ,
    \msto[13][hwrite] ,
    \msto[13][hsize] ,
    \msto[13][hburst] ,
    \msto[13][hprot] ,
    \msto[13][hwdata] ,
    \msto[13][hirq] ,
    \msto[13][hconfig][0] ,
    \msto[13][hconfig][1] ,
    \msto[13][hconfig][2] ,
    \msto[13][hconfig][3] ,
    \msto[13][hconfig][4] ,
    \msto[13][hconfig][5] ,
    \msto[13][hconfig][6] ,
    \msto[13][hconfig][7] ,
    \msto[13][hindex] ,
    \msto[12][hbusreq] ,
    \msto[12][hlock] ,
    \msto[12][htrans] ,
    \msto[12][haddr] ,
    \msto[12][hwrite] ,
    \msto[12][hsize] ,
    \msto[12][hburst] ,
    \msto[12][hprot] ,
    \msto[12][hwdata] ,
    \msto[12][hirq] ,
    \msto[12][hconfig][0] ,
    \msto[12][hconfig][1] ,
    \msto[12][hconfig][2] ,
    \msto[12][hconfig][3] ,
    \msto[12][hconfig][4] ,
    \msto[12][hconfig][5] ,
    \msto[12][hconfig][6] ,
    \msto[12][hconfig][7] ,
    \msto[12][hindex] ,
    \msto[11][hbusreq] ,
    \msto[11][hlock] ,
    \msto[11][htrans] ,
    \msto[11][haddr] ,
    \msto[11][hwrite] ,
    \msto[11][hsize] ,
    \msto[11][hburst] ,
    \msto[11][hprot] ,
    \msto[11][hwdata] ,
    \msto[11][hirq] ,
    \msto[11][hconfig][0] ,
    \msto[11][hconfig][1] ,
    \msto[11][hconfig][2] ,
    \msto[11][hconfig][3] ,
    \msto[11][hconfig][4] ,
    \msto[11][hconfig][5] ,
    \msto[11][hconfig][6] ,
    \msto[11][hconfig][7] ,
    \msto[11][hindex] ,
    \msto[10][hbusreq] ,
    \msto[10][hlock] ,
    \msto[10][htrans] ,
    \msto[10][haddr] ,
    \msto[10][hwrite] ,
    \msto[10][hsize] ,
    \msto[10][hburst] ,
    \msto[10][hprot] ,
    \msto[10][hwdata] ,
    \msto[10][hirq] ,
    \msto[10][hconfig][0] ,
    \msto[10][hconfig][1] ,
    \msto[10][hconfig][2] ,
    \msto[10][hconfig][3] ,
    \msto[10][hconfig][4] ,
    \msto[10][hconfig][5] ,
    \msto[10][hconfig][6] ,
    \msto[10][hconfig][7] ,
    \msto[10][hindex] ,
    \msto[9][hbusreq] ,
    \msto[9][hlock] ,
    \msto[9][htrans] ,
    \msto[9][haddr] ,
    \msto[9][hwrite] ,
    \msto[9][hsize] ,
    \msto[9][hburst] ,
    \msto[9][hprot] ,
    \msto[9][hwdata] ,
    \msto[9][hirq] ,
    \msto[9][hconfig][0] ,
    \msto[9][hconfig][1] ,
    \msto[9][hconfig][2] ,
    \msto[9][hconfig][3] ,
    \msto[9][hconfig][4] ,
    \msto[9][hconfig][5] ,
    \msto[9][hconfig][6] ,
    \msto[9][hconfig][7] ,
    \msto[9][hindex] ,
    \msto[8][hbusreq] ,
    \msto[8][hlock] ,
    \msto[8][htrans] ,
    \msto[8][haddr] ,
    \msto[8][hwrite] ,
    \msto[8][hsize] ,
    \msto[8][hburst] ,
    \msto[8][hprot] ,
    \msto[8][hwdata] ,
    \msto[8][hirq] ,
    \msto[8][hconfig][0] ,
    \msto[8][hconfig][1] ,
    \msto[8][hconfig][2] ,
    \msto[8][hconfig][3] ,
    \msto[8][hconfig][4] ,
    \msto[8][hconfig][5] ,
    \msto[8][hconfig][6] ,
    \msto[8][hconfig][7] ,
    \msto[8][hindex] ,
    .\msto[7][hbusreq] (msto),
    \msto[7][hlock] ,
    \msto[7][htrans] ,
    \msto[7][haddr] ,
    \msto[7][hwrite] ,
    \msto[7][hsize] ,
    \msto[7][hburst] ,
    \msto[7][hprot] ,
    \msto[7][hwdata] ,
    \msto[7][hirq] ,
    \msto[7][hconfig][0] ,
    \msto[7][hconfig][1] ,
    \msto[7][hconfig][2] ,
    \msto[7][hconfig][3] ,
    \msto[7][hconfig][4] ,
    \msto[7][hconfig][5] ,
    \msto[7][hconfig][6] ,
    \msto[7][hconfig][7] ,
    \msto[7][hindex] ,
    \msto[6][hbusreq] ,
    \msto[6][hlock] ,
    \msto[6][htrans] ,
    \msto[6][haddr] ,
    \msto[6][hwrite] ,
    \msto[6][hsize] ,
    \msto[6][hburst] ,
    \msto[6][hprot] ,
    \msto[6][hwdata] ,
    \msto[6][hirq] ,
    \msto[6][hconfig][0] ,
    \msto[6][hconfig][1] ,
    \msto[6][hconfig][2] ,
    \msto[6][hconfig][3] ,
    \msto[6][hconfig][4] ,
    \msto[6][hconfig][5] ,
    \msto[6][hconfig][6] ,
    \msto[6][hconfig][7] ,
    \msto[6][hindex] ,
    \msto[5][hbusreq] ,
    \msto[5][hlock] ,
    \msto[5][htrans] ,
    \msto[5][haddr] ,
    \msto[5][hwrite] ,
    \msto[5][hsize] ,
    \msto[5][hburst] ,
    \msto[5][hprot] ,
    \msto[5][hwdata] ,
    \msto[5][hirq] ,
    \msto[5][hconfig][0] ,
    \msto[5][hconfig][1] ,
    \msto[5][hconfig][2] ,
    \msto[5][hconfig][3] ,
    \msto[5][hconfig][4] ,
    \msto[5][hconfig][5] ,
    \msto[5][hconfig][6] ,
    \msto[5][hconfig][7] ,
    \msto[5][hindex] ,
    \msto[4][hbusreq] ,
    \msto[4][hlock] ,
    \msto[4][htrans] ,
    \msto[4][haddr] ,
    \msto[4][hwrite] ,
    \msto[4][hsize] ,
    \msto[4][hburst] ,
    \msto[4][hprot] ,
    \msto[4][hwdata] ,
    \msto[4][hirq] ,
    \msto[4][hconfig][0] ,
    \msto[4][hconfig][1] ,
    \msto[4][hconfig][2] ,
    \msto[4][hconfig][3] ,
    \msto[4][hconfig][4] ,
    \msto[4][hconfig][5] ,
    \msto[4][hconfig][6] ,
    \msto[4][hconfig][7] ,
    \msto[4][hindex] ,
    \msto[3][hbusreq] ,
    \msto[3][hlock] ,
    \msto[3][htrans] ,
    \msto[3][haddr] ,
    \msto[3][hwrite] ,
    \msto[3][hsize] ,
    \msto[3][hburst] ,
    \msto[3][hprot] ,
    \msto[3][hwdata] ,
    \msto[3][hirq] ,
    \msto[3][hconfig][0] ,
    \msto[3][hconfig][1] ,
    \msto[3][hconfig][2] ,
    \msto[3][hconfig][3] ,
    \msto[3][hconfig][4] ,
    \msto[3][hconfig][5] ,
    \msto[3][hconfig][6] ,
    \msto[3][hconfig][7] ,
    \msto[3][hindex] ,
    \msto[2][hbusreq] ,
    \msto[2][hlock] ,
    \msto[2][htrans] ,
    \msto[2][haddr] ,
    \msto[2][hwrite] ,
    \msto[2][hsize] ,
    \msto[2][hburst] ,
    \msto[2][hprot] ,
    \msto[2][hwdata] ,
    \msto[2][hirq] ,
    \msto[2][hconfig][0] ,
    \msto[2][hconfig][1] ,
    \msto[2][hconfig][2] ,
    \msto[2][hconfig][3] ,
    \msto[2][hconfig][4] ,
    \msto[2][hconfig][5] ,
    \msto[2][hconfig][6] ,
    \msto[2][hconfig][7] ,
    \msto[2][hindex] ,
    \msto[1][hbusreq] ,
    \msto[1][hlock] ,
    \msto[1][htrans] ,
    \msto[1][haddr] ,
    \msto[1][hwrite] ,
    \msto[1][hsize] ,
    \msto[1][hburst] ,
    \msto[1][hprot] ,
    \msto[1][hwdata] ,
    \msto[1][hirq] ,
    \msto[1][hconfig][0] ,
    \msto[1][hconfig][1] ,
    \msto[1][hconfig][2] ,
    \msto[1][hconfig][3] ,
    \msto[1][hconfig][4] ,
    \msto[1][hconfig][5] ,
    \msto[1][hconfig][6] ,
    \msto[1][hconfig][7] ,
    \msto[1][hindex] ,
    \msto[0][hbusreq] ,
    \msto[0][hlock] ,
    \msto[0][htrans] ,
    \msto[0][haddr] ,
    \msto[0][hwrite] ,
    \msto[0][hsize] ,
    \msto[0][hburst] ,
    \msto[0][hprot] ,
    \msto[0][hwdata] ,
    \msto[0][hirq] ,
    \msto[0][hconfig][0] ,
    \msto[0][hconfig][1] ,
    \msto[0][hconfig][2] ,
    \msto[0][hconfig][3] ,
    \msto[0][hconfig][4] ,
    \msto[0][hconfig][5] ,
    \msto[0][hconfig][6] ,
    \msto[0][hconfig][7] ,
    \msto[0][hindex] ,
    \slvi[hsel] ,
    \slvi[haddr] ,
    \slvi[hwrite] ,
    \slvi[htrans] ,
    \slvi[hsize] ,
    \slvi[hburst] ,
    \slvi[hwdata] ,
    \slvi[hprot] ,
    \slvi[hready] ,
    \slvi[hmaster] ,
    \slvi[hmastlock] ,
    \slvi[hmbsel] ,
    \slvi[hirq] ,
    \slvi[testen] ,
    \slvi[testrst] ,
    \slvi[scanen] ,
    \slvi[testoen] ,
    \slvi[testin] ,
    \slvo[15][hready] ,
    \slvo[15][hresp] ,
    \slvo[15][hrdata] ,
    \slvo[15][hsplit] ,
    \slvo[15][hirq] ,
    \slvo[15][hconfig][0] ,
    \slvo[15][hconfig][1] ,
    \slvo[15][hconfig][2] ,
    \slvo[15][hconfig][3] ,
    \slvo[15][hconfig][4] ,
    \slvo[15][hconfig][5] ,
    \slvo[15][hconfig][6] ,
    \slvo[15][hconfig][7] ,
    \slvo[15][hindex] ,
    \slvo[14][hready] ,
    \slvo[14][hresp] ,
    \slvo[14][hrdata] ,
    \slvo[14][hsplit] ,
    \slvo[14][hirq] ,
    \slvo[14][hconfig][0] ,
    \slvo[14][hconfig][1] ,
    \slvo[14][hconfig][2] ,
    \slvo[14][hconfig][3] ,
    \slvo[14][hconfig][4] ,
    \slvo[14][hconfig][5] ,
    \slvo[14][hconfig][6] ,
    \slvo[14][hconfig][7] ,
    \slvo[14][hindex] ,
    \slvo[13][hready] ,
    \slvo[13][hresp] ,
    \slvo[13][hrdata] ,
    \slvo[13][hsplit] ,
    \slvo[13][hirq] ,
    \slvo[13][hconfig][0] ,
    \slvo[13][hconfig][1] ,
    \slvo[13][hconfig][2] ,
    \slvo[13][hconfig][3] ,
    \slvo[13][hconfig][4] ,
    \slvo[13][hconfig][5] ,
    \slvo[13][hconfig][6] ,
    \slvo[13][hconfig][7] ,
    \slvo[13][hindex] ,
    \slvo[12][hready] ,
    \slvo[12][hresp] ,
    \slvo[12][hrdata] ,
    \slvo[12][hsplit] ,
    \slvo[12][hirq] ,
    \slvo[12][hconfig][0] ,
    \slvo[12][hconfig][1] ,
    \slvo[12][hconfig][2] ,
    \slvo[12][hconfig][3] ,
    \slvo[12][hconfig][4] ,
    \slvo[12][hconfig][5] ,
    \slvo[12][hconfig][6] ,
    \slvo[12][hconfig][7] ,
    \slvo[12][hindex] ,
    \slvo[11][hready] ,
    \slvo[11][hresp] ,
    \slvo[11][hrdata] ,
    \slvo[11][hsplit] ,
    \slvo[11][hirq] ,
    \slvo[11][hconfig][0] ,
    \slvo[11][hconfig][1] ,
    \slvo[11][hconfig][2] ,
    \slvo[11][hconfig][3] ,
    \slvo[11][hconfig][4] ,
    \slvo[11][hconfig][5] ,
    \slvo[11][hconfig][6] ,
    \slvo[11][hconfig][7] ,
    \slvo[11][hindex] ,
    \slvo[10][hready] ,
    \slvo[10][hresp] ,
    \slvo[10][hrdata] ,
    \slvo[10][hsplit] ,
    \slvo[10][hirq] ,
    \slvo[10][hconfig][0] ,
    \slvo[10][hconfig][1] ,
    \slvo[10][hconfig][2] ,
    \slvo[10][hconfig][3] ,
    \slvo[10][hconfig][4] ,
    \slvo[10][hconfig][5] ,
    \slvo[10][hconfig][6] ,
    \slvo[10][hconfig][7] ,
    \slvo[10][hindex] ,
    \slvo[9][hready] ,
    \slvo[9][hresp] ,
    \slvo[9][hrdata] ,
    \slvo[9][hsplit] ,
    \slvo[9][hirq] ,
    \slvo[9][hconfig][0] ,
    \slvo[9][hconfig][1] ,
    \slvo[9][hconfig][2] ,
    \slvo[9][hconfig][3] ,
    \slvo[9][hconfig][4] ,
    \slvo[9][hconfig][5] ,
    \slvo[9][hconfig][6] ,
    \slvo[9][hconfig][7] ,
    \slvo[9][hindex] ,
    \slvo[8][hready] ,
    \slvo[8][hresp] ,
    \slvo[8][hrdata] ,
    \slvo[8][hsplit] ,
    \slvo[8][hirq] ,
    \slvo[8][hconfig][0] ,
    \slvo[8][hconfig][1] ,
    \slvo[8][hconfig][2] ,
    \slvo[8][hconfig][3] ,
    \slvo[8][hconfig][4] ,
    \slvo[8][hconfig][5] ,
    \slvo[8][hconfig][6] ,
    \slvo[8][hconfig][7] ,
    \slvo[8][hindex] ,
    .\slvo[7][hready] (slvo),
    \slvo[7][hresp] ,
    \slvo[7][hrdata] ,
    \slvo[7][hsplit] ,
    \slvo[7][hirq] ,
    \slvo[7][hconfig][0] ,
    \slvo[7][hconfig][1] ,
    \slvo[7][hconfig][2] ,
    \slvo[7][hconfig][3] ,
    \slvo[7][hconfig][4] ,
    \slvo[7][hconfig][5] ,
    \slvo[7][hconfig][6] ,
    \slvo[7][hconfig][7] ,
    \slvo[7][hindex] ,
    \slvo[6][hready] ,
    \slvo[6][hresp] ,
    \slvo[6][hrdata] ,
    \slvo[6][hsplit] ,
    \slvo[6][hirq] ,
    \slvo[6][hconfig][0] ,
    \slvo[6][hconfig][1] ,
    \slvo[6][hconfig][2] ,
    \slvo[6][hconfig][3] ,
    \slvo[6][hconfig][4] ,
    \slvo[6][hconfig][5] ,
    \slvo[6][hconfig][6] ,
    \slvo[6][hconfig][7] ,
    \slvo[6][hindex] ,
    \slvo[5][hready] ,
    \slvo[5][hresp] ,
    \slvo[5][hrdata] ,
    \slvo[5][hsplit] ,
    \slvo[5][hirq] ,
    \slvo[5][hconfig][0] ,
    \slvo[5][hconfig][1] ,
    \slvo[5][hconfig][2] ,
    \slvo[5][hconfig][3] ,
    \slvo[5][hconfig][4] ,
    \slvo[5][hconfig][5] ,
    \slvo[5][hconfig][6] ,
    \slvo[5][hconfig][7] ,
    \slvo[5][hindex] ,
    \slvo[4][hready] ,
    \slvo[4][hresp] ,
    \slvo[4][hrdata] ,
    \slvo[4][hsplit] ,
    \slvo[4][hirq] ,
    \slvo[4][hconfig][0] ,
    \slvo[4][hconfig][1] ,
    \slvo[4][hconfig][2] ,
    \slvo[4][hconfig][3] ,
    \slvo[4][hconfig][4] ,
    \slvo[4][hconfig][5] ,
    \slvo[4][hconfig][6] ,
    \slvo[4][hconfig][7] ,
    \slvo[4][hindex] ,
    \slvo[3][hready] ,
    \slvo[3][hresp] ,
    \slvo[3][hrdata] ,
    \slvo[3][hsplit] ,
    \slvo[3][hirq] ,
    \slvo[3][hconfig][0] ,
    \slvo[3][hconfig][1] ,
    \slvo[3][hconfig][2] ,
    \slvo[3][hconfig][3] ,
    \slvo[3][hconfig][4] ,
    \slvo[3][hconfig][5] ,
    \slvo[3][hconfig][6] ,
    \slvo[3][hconfig][7] ,
    \slvo[3][hindex] ,
    \slvo[2][hready] ,
    \slvo[2][hresp] ,
    \slvo[2][hrdata] ,
    \slvo[2][hsplit] ,
    \slvo[2][hirq] ,
    \slvo[2][hconfig][0] ,
    \slvo[2][hconfig][1] ,
    \slvo[2][hconfig][2] ,
    \slvo[2][hconfig][3] ,
    \slvo[2][hconfig][4] ,
    \slvo[2][hconfig][5] ,
    \slvo[2][hconfig][6] ,
    \slvo[2][hconfig][7] ,
    \slvo[2][hindex] ,
    \slvo[1][hready] ,
    \slvo[1][hresp] ,
    \slvo[1][hrdata] ,
    \slvo[1][hsplit] ,
    \slvo[1][hirq] ,
    \slvo[1][hconfig][0] ,
    \slvo[1][hconfig][1] ,
    \slvo[1][hconfig][2] ,
    \slvo[1][hconfig][3] ,
    \slvo[1][hconfig][4] ,
    \slvo[1][hconfig][5] ,
    \slvo[1][hconfig][6] ,
    \slvo[1][hconfig][7] ,
    \slvo[1][hindex] ,
    \slvo[0][hready] ,
    \slvo[0][hresp] ,
    \slvo[0][hrdata] ,
    \slvo[0][hsplit] ,
    \slvo[0][hirq] ,
    \slvo[0][hconfig][0] ,
    \slvo[0][hconfig][1] ,
    \slvo[0][hconfig][2] ,
    \slvo[0][hconfig][3] ,
    \slvo[0][hconfig][4] ,
    \slvo[0][hconfig][5] ,
    \slvo[0][hconfig][6] ,
    \slvo[0][hconfig][7] ,
    \slvo[0][hindex] ,
    testen,
    testrst,
    scanen,
    testoen,
    testsig);
  input rst;
  input clk;
  output [0:15]\msti[hgrant] ;
  output \msti[hready] ;
  output [1:0]\msti[hresp] ;
  output [31:0]\msti[hrdata] ;
  output [31:0]\msti[hirq] ;
  output \msti[testen] ;
  output \msti[testrst] ;
  output \msti[scanen] ;
  output \msti[testoen] ;
  output [3:0]\msti[testin] ;
  input \msto[15][hbusreq] ;
  input \msto[15][hlock] ;
  input [1:0]\msto[15][htrans] ;
  input [31:0]\msto[15][haddr] ;
  input \msto[15][hwrite] ;
  input [2:0]\msto[15][hsize] ;
  input [2:0]\msto[15][hburst] ;
  input [3:0]\msto[15][hprot] ;
  input [31:0]\msto[15][hwdata] ;
  input [31:0]\msto[15][hirq] ;
  input [31:0]\msto[15][hconfig][0] ;
  input [31:0]\msto[15][hconfig][1] ;
  input [31:0]\msto[15][hconfig][2] ;
  input [31:0]\msto[15][hconfig][3] ;
  input [31:0]\msto[15][hconfig][4] ;
  input [31:0]\msto[15][hconfig][5] ;
  input [31:0]\msto[15][hconfig][6] ;
  input [31:0]\msto[15][hconfig][7] ;
  input [3:0]\msto[15][hindex] ;
  input \msto[14][hbusreq] ;
  input \msto[14][hlock] ;
  input [1:0]\msto[14][htrans] ;
  input [31:0]\msto[14][haddr] ;
  input \msto[14][hwrite] ;
  input [2:0]\msto[14][hsize] ;
  input [2:0]\msto[14][hburst] ;
  input [3:0]\msto[14][hprot] ;
  input [31:0]\msto[14][hwdata] ;
  input [31:0]\msto[14][hirq] ;
  input [31:0]\msto[14][hconfig][0] ;
  input [31:0]\msto[14][hconfig][1] ;
  input [31:0]\msto[14][hconfig][2] ;
  input [31:0]\msto[14][hconfig][3] ;
  input [31:0]\msto[14][hconfig][4] ;
  input [31:0]\msto[14][hconfig][5] ;
  input [31:0]\msto[14][hconfig][6] ;
  input [31:0]\msto[14][hconfig][7] ;
  input [3:0]\msto[14][hindex] ;
  input \msto[13][hbusreq] ;
  input \msto[13][hlock] ;
  input [1:0]\msto[13][htrans] ;
  input [31:0]\msto[13][haddr] ;
  input \msto[13][hwrite] ;
  input [2:0]\msto[13][hsize] ;
  input [2:0]\msto[13][hburst] ;
  input [3:0]\msto[13][hprot] ;
  input [31:0]\msto[13][hwdata] ;
  input [31:0]\msto[13][hirq] ;
  input [31:0]\msto[13][hconfig][0] ;
  input [31:0]\msto[13][hconfig][1] ;
  input [31:0]\msto[13][hconfig][2] ;
  input [31:0]\msto[13][hconfig][3] ;
  input [31:0]\msto[13][hconfig][4] ;
  input [31:0]\msto[13][hconfig][5] ;
  input [31:0]\msto[13][hconfig][6] ;
  input [31:0]\msto[13][hconfig][7] ;
  input [3:0]\msto[13][hindex] ;
  input \msto[12][hbusreq] ;
  input \msto[12][hlock] ;
  input [1:0]\msto[12][htrans] ;
  input [31:0]\msto[12][haddr] ;
  input \msto[12][hwrite] ;
  input [2:0]\msto[12][hsize] ;
  input [2:0]\msto[12][hburst] ;
  input [3:0]\msto[12][hprot] ;
  input [31:0]\msto[12][hwdata] ;
  input [31:0]\msto[12][hirq] ;
  input [31:0]\msto[12][hconfig][0] ;
  input [31:0]\msto[12][hconfig][1] ;
  input [31:0]\msto[12][hconfig][2] ;
  input [31:0]\msto[12][hconfig][3] ;
  input [31:0]\msto[12][hconfig][4] ;
  input [31:0]\msto[12][hconfig][5] ;
  input [31:0]\msto[12][hconfig][6] ;
  input [31:0]\msto[12][hconfig][7] ;
  input [3:0]\msto[12][hindex] ;
  input \msto[11][hbusreq] ;
  input \msto[11][hlock] ;
  input [1:0]\msto[11][htrans] ;
  input [31:0]\msto[11][haddr] ;
  input \msto[11][hwrite] ;
  input [2:0]\msto[11][hsize] ;
  input [2:0]\msto[11][hburst] ;
  input [3:0]\msto[11][hprot] ;
  input [31:0]\msto[11][hwdata] ;
  input [31:0]\msto[11][hirq] ;
  input [31:0]\msto[11][hconfig][0] ;
  input [31:0]\msto[11][hconfig][1] ;
  input [31:0]\msto[11][hconfig][2] ;
  input [31:0]\msto[11][hconfig][3] ;
  input [31:0]\msto[11][hconfig][4] ;
  input [31:0]\msto[11][hconfig][5] ;
  input [31:0]\msto[11][hconfig][6] ;
  input [31:0]\msto[11][hconfig][7] ;
  input [3:0]\msto[11][hindex] ;
  input \msto[10][hbusreq] ;
  input \msto[10][hlock] ;
  input [1:0]\msto[10][htrans] ;
  input [31:0]\msto[10][haddr] ;
  input \msto[10][hwrite] ;
  input [2:0]\msto[10][hsize] ;
  input [2:0]\msto[10][hburst] ;
  input [3:0]\msto[10][hprot] ;
  input [31:0]\msto[10][hwdata] ;
  input [31:0]\msto[10][hirq] ;
  input [31:0]\msto[10][hconfig][0] ;
  input [31:0]\msto[10][hconfig][1] ;
  input [31:0]\msto[10][hconfig][2] ;
  input [31:0]\msto[10][hconfig][3] ;
  input [31:0]\msto[10][hconfig][4] ;
  input [31:0]\msto[10][hconfig][5] ;
  input [31:0]\msto[10][hconfig][6] ;
  input [31:0]\msto[10][hconfig][7] ;
  input [3:0]\msto[10][hindex] ;
  input \msto[9][hbusreq] ;
  input \msto[9][hlock] ;
  input [1:0]\msto[9][htrans] ;
  input [31:0]\msto[9][haddr] ;
  input \msto[9][hwrite] ;
  input [2:0]\msto[9][hsize] ;
  input [2:0]\msto[9][hburst] ;
  input [3:0]\msto[9][hprot] ;
  input [31:0]\msto[9][hwdata] ;
  input [31:0]\msto[9][hirq] ;
  input [31:0]\msto[9][hconfig][0] ;
  input [31:0]\msto[9][hconfig][1] ;
  input [31:0]\msto[9][hconfig][2] ;
  input [31:0]\msto[9][hconfig][3] ;
  input [31:0]\msto[9][hconfig][4] ;
  input [31:0]\msto[9][hconfig][5] ;
  input [31:0]\msto[9][hconfig][6] ;
  input [31:0]\msto[9][hconfig][7] ;
  input [3:0]\msto[9][hindex] ;
  input \msto[8][hbusreq] ;
  input \msto[8][hlock] ;
  input [1:0]\msto[8][htrans] ;
  input [31:0]\msto[8][haddr] ;
  input \msto[8][hwrite] ;
  input [2:0]\msto[8][hsize] ;
  input [2:0]\msto[8][hburst] ;
  input [3:0]\msto[8][hprot] ;
  input [31:0]\msto[8][hwdata] ;
  input [31:0]\msto[8][hirq] ;
  input [31:0]\msto[8][hconfig][0] ;
  input [31:0]\msto[8][hconfig][1] ;
  input [31:0]\msto[8][hconfig][2] ;
  input [31:0]\msto[8][hconfig][3] ;
  input [31:0]\msto[8][hconfig][4] ;
  input [31:0]\msto[8][hconfig][5] ;
  input [31:0]\msto[8][hconfig][6] ;
  input [31:0]\msto[8][hconfig][7] ;
  input [3:0]\msto[8][hindex] ;
  input \msto[7][hlock] ;
  input [1:0]\msto[7][htrans] ;
  input [31:0]\msto[7][haddr] ;
  input \msto[7][hwrite] ;
  input [2:0]\msto[7][hsize] ;
  input [2:0]\msto[7][hburst] ;
  input [3:0]\msto[7][hprot] ;
  input [31:0]\msto[7][hwdata] ;
  input [31:0]\msto[7][hirq] ;
  input [31:0]\msto[7][hconfig][0] ;
  input [31:0]\msto[7][hconfig][1] ;
  input [31:0]\msto[7][hconfig][2] ;
  input [31:0]\msto[7][hconfig][3] ;
  input [31:0]\msto[7][hconfig][4] ;
  input [31:0]\msto[7][hconfig][5] ;
  input [31:0]\msto[7][hconfig][6] ;
  input [31:0]\msto[7][hconfig][7] ;
  input [3:0]\msto[7][hindex] ;
  input \msto[6][hbusreq] ;
  input \msto[6][hlock] ;
  input [1:0]\msto[6][htrans] ;
  input [31:0]\msto[6][haddr] ;
  input \msto[6][hwrite] ;
  input [2:0]\msto[6][hsize] ;
  input [2:0]\msto[6][hburst] ;
  input [3:0]\msto[6][hprot] ;
  input [31:0]\msto[6][hwdata] ;
  input [31:0]\msto[6][hirq] ;
  input [31:0]\msto[6][hconfig][0] ;
  input [31:0]\msto[6][hconfig][1] ;
  input [31:0]\msto[6][hconfig][2] ;
  input [31:0]\msto[6][hconfig][3] ;
  input [31:0]\msto[6][hconfig][4] ;
  input [31:0]\msto[6][hconfig][5] ;
  input [31:0]\msto[6][hconfig][6] ;
  input [31:0]\msto[6][hconfig][7] ;
  input [3:0]\msto[6][hindex] ;
  input \msto[5][hbusreq] ;
  input \msto[5][hlock] ;
  input [1:0]\msto[5][htrans] ;
  input [31:0]\msto[5][haddr] ;
  input \msto[5][hwrite] ;
  input [2:0]\msto[5][hsize] ;
  input [2:0]\msto[5][hburst] ;
  input [3:0]\msto[5][hprot] ;
  input [31:0]\msto[5][hwdata] ;
  input [31:0]\msto[5][hirq] ;
  input [31:0]\msto[5][hconfig][0] ;
  input [31:0]\msto[5][hconfig][1] ;
  input [31:0]\msto[5][hconfig][2] ;
  input [31:0]\msto[5][hconfig][3] ;
  input [31:0]\msto[5][hconfig][4] ;
  input [31:0]\msto[5][hconfig][5] ;
  input [31:0]\msto[5][hconfig][6] ;
  input [31:0]\msto[5][hconfig][7] ;
  input [3:0]\msto[5][hindex] ;
  input \msto[4][hbusreq] ;
  input \msto[4][hlock] ;
  input [1:0]\msto[4][htrans] ;
  input [31:0]\msto[4][haddr] ;
  input \msto[4][hwrite] ;
  input [2:0]\msto[4][hsize] ;
  input [2:0]\msto[4][hburst] ;
  input [3:0]\msto[4][hprot] ;
  input [31:0]\msto[4][hwdata] ;
  input [31:0]\msto[4][hirq] ;
  input [31:0]\msto[4][hconfig][0] ;
  input [31:0]\msto[4][hconfig][1] ;
  input [31:0]\msto[4][hconfig][2] ;
  input [31:0]\msto[4][hconfig][3] ;
  input [31:0]\msto[4][hconfig][4] ;
  input [31:0]\msto[4][hconfig][5] ;
  input [31:0]\msto[4][hconfig][6] ;
  input [31:0]\msto[4][hconfig][7] ;
  input [3:0]\msto[4][hindex] ;
  input \msto[3][hbusreq] ;
  input \msto[3][hlock] ;
  input [1:0]\msto[3][htrans] ;
  input [31:0]\msto[3][haddr] ;
  input \msto[3][hwrite] ;
  input [2:0]\msto[3][hsize] ;
  input [2:0]\msto[3][hburst] ;
  input [3:0]\msto[3][hprot] ;
  input [31:0]\msto[3][hwdata] ;
  input [31:0]\msto[3][hirq] ;
  input [31:0]\msto[3][hconfig][0] ;
  input [31:0]\msto[3][hconfig][1] ;
  input [31:0]\msto[3][hconfig][2] ;
  input [31:0]\msto[3][hconfig][3] ;
  input [31:0]\msto[3][hconfig][4] ;
  input [31:0]\msto[3][hconfig][5] ;
  input [31:0]\msto[3][hconfig][6] ;
  input [31:0]\msto[3][hconfig][7] ;
  input [3:0]\msto[3][hindex] ;
  input \msto[2][hbusreq] ;
  input \msto[2][hlock] ;
  input [1:0]\msto[2][htrans] ;
  input [31:0]\msto[2][haddr] ;
  input \msto[2][hwrite] ;
  input [2:0]\msto[2][hsize] ;
  input [2:0]\msto[2][hburst] ;
  input [3:0]\msto[2][hprot] ;
  input [31:0]\msto[2][hwdata] ;
  input [31:0]\msto[2][hirq] ;
  input [31:0]\msto[2][hconfig][0] ;
  input [31:0]\msto[2][hconfig][1] ;
  input [31:0]\msto[2][hconfig][2] ;
  input [31:0]\msto[2][hconfig][3] ;
  input [31:0]\msto[2][hconfig][4] ;
  input [31:0]\msto[2][hconfig][5] ;
  input [31:0]\msto[2][hconfig][6] ;
  input [31:0]\msto[2][hconfig][7] ;
  input [3:0]\msto[2][hindex] ;
  input \msto[1][hbusreq] ;
  input \msto[1][hlock] ;
  input [1:0]\msto[1][htrans] ;
  input [31:0]\msto[1][haddr] ;
  input \msto[1][hwrite] ;
  input [2:0]\msto[1][hsize] ;
  input [2:0]\msto[1][hburst] ;
  input [3:0]\msto[1][hprot] ;
  input [31:0]\msto[1][hwdata] ;
  input [31:0]\msto[1][hirq] ;
  input [31:0]\msto[1][hconfig][0] ;
  input [31:0]\msto[1][hconfig][1] ;
  input [31:0]\msto[1][hconfig][2] ;
  input [31:0]\msto[1][hconfig][3] ;
  input [31:0]\msto[1][hconfig][4] ;
  input [31:0]\msto[1][hconfig][5] ;
  input [31:0]\msto[1][hconfig][6] ;
  input [31:0]\msto[1][hconfig][7] ;
  input [3:0]\msto[1][hindex] ;
  input \msto[0][hbusreq] ;
  input \msto[0][hlock] ;
  input [1:0]\msto[0][htrans] ;
  input [31:0]\msto[0][haddr] ;
  input \msto[0][hwrite] ;
  input [2:0]\msto[0][hsize] ;
  input [2:0]\msto[0][hburst] ;
  input [3:0]\msto[0][hprot] ;
  input [31:0]\msto[0][hwdata] ;
  input [31:0]\msto[0][hirq] ;
  input [31:0]\msto[0][hconfig][0] ;
  input [31:0]\msto[0][hconfig][1] ;
  input [31:0]\msto[0][hconfig][2] ;
  input [31:0]\msto[0][hconfig][3] ;
  input [31:0]\msto[0][hconfig][4] ;
  input [31:0]\msto[0][hconfig][5] ;
  input [31:0]\msto[0][hconfig][6] ;
  input [31:0]\msto[0][hconfig][7] ;
  input [3:0]\msto[0][hindex] ;
  output [0:15]\slvi[hsel] ;
  output [31:0]\slvi[haddr] ;
  output \slvi[hwrite] ;
  output [1:0]\slvi[htrans] ;
  output [2:0]\slvi[hsize] ;
  output [2:0]\slvi[hburst] ;
  output [31:0]\slvi[hwdata] ;
  output [3:0]\slvi[hprot] ;
  output \slvi[hready] ;
  output [3:0]\slvi[hmaster] ;
  output \slvi[hmastlock] ;
  output [0:3]\slvi[hmbsel] ;
  output [31:0]\slvi[hirq] ;
  output \slvi[testen] ;
  output \slvi[testrst] ;
  output \slvi[scanen] ;
  output \slvi[testoen] ;
  output [3:0]\slvi[testin] ;
  input \slvo[15][hready] ;
  input [1:0]\slvo[15][hresp] ;
  input [31:0]\slvo[15][hrdata] ;
  input [15:0]\slvo[15][hsplit] ;
  input [31:0]\slvo[15][hirq] ;
  input [31:0]\slvo[15][hconfig][0] ;
  input [31:0]\slvo[15][hconfig][1] ;
  input [31:0]\slvo[15][hconfig][2] ;
  input [31:0]\slvo[15][hconfig][3] ;
  input [31:0]\slvo[15][hconfig][4] ;
  input [31:0]\slvo[15][hconfig][5] ;
  input [31:0]\slvo[15][hconfig][6] ;
  input [31:0]\slvo[15][hconfig][7] ;
  input [3:0]\slvo[15][hindex] ;
  input \slvo[14][hready] ;
  input [1:0]\slvo[14][hresp] ;
  input [31:0]\slvo[14][hrdata] ;
  input [15:0]\slvo[14][hsplit] ;
  input [31:0]\slvo[14][hirq] ;
  input [31:0]\slvo[14][hconfig][0] ;
  input [31:0]\slvo[14][hconfig][1] ;
  input [31:0]\slvo[14][hconfig][2] ;
  input [31:0]\slvo[14][hconfig][3] ;
  input [31:0]\slvo[14][hconfig][4] ;
  input [31:0]\slvo[14][hconfig][5] ;
  input [31:0]\slvo[14][hconfig][6] ;
  input [31:0]\slvo[14][hconfig][7] ;
  input [3:0]\slvo[14][hindex] ;
  input \slvo[13][hready] ;
  input [1:0]\slvo[13][hresp] ;
  input [31:0]\slvo[13][hrdata] ;
  input [15:0]\slvo[13][hsplit] ;
  input [31:0]\slvo[13][hirq] ;
  input [31:0]\slvo[13][hconfig][0] ;
  input [31:0]\slvo[13][hconfig][1] ;
  input [31:0]\slvo[13][hconfig][2] ;
  input [31:0]\slvo[13][hconfig][3] ;
  input [31:0]\slvo[13][hconfig][4] ;
  input [31:0]\slvo[13][hconfig][5] ;
  input [31:0]\slvo[13][hconfig][6] ;
  input [31:0]\slvo[13][hconfig][7] ;
  input [3:0]\slvo[13][hindex] ;
  input \slvo[12][hready] ;
  input [1:0]\slvo[12][hresp] ;
  input [31:0]\slvo[12][hrdata] ;
  input [15:0]\slvo[12][hsplit] ;
  input [31:0]\slvo[12][hirq] ;
  input [31:0]\slvo[12][hconfig][0] ;
  input [31:0]\slvo[12][hconfig][1] ;
  input [31:0]\slvo[12][hconfig][2] ;
  input [31:0]\slvo[12][hconfig][3] ;
  input [31:0]\slvo[12][hconfig][4] ;
  input [31:0]\slvo[12][hconfig][5] ;
  input [31:0]\slvo[12][hconfig][6] ;
  input [31:0]\slvo[12][hconfig][7] ;
  input [3:0]\slvo[12][hindex] ;
  input \slvo[11][hready] ;
  input [1:0]\slvo[11][hresp] ;
  input [31:0]\slvo[11][hrdata] ;
  input [15:0]\slvo[11][hsplit] ;
  input [31:0]\slvo[11][hirq] ;
  input [31:0]\slvo[11][hconfig][0] ;
  input [31:0]\slvo[11][hconfig][1] ;
  input [31:0]\slvo[11][hconfig][2] ;
  input [31:0]\slvo[11][hconfig][3] ;
  input [31:0]\slvo[11][hconfig][4] ;
  input [31:0]\slvo[11][hconfig][5] ;
  input [31:0]\slvo[11][hconfig][6] ;
  input [31:0]\slvo[11][hconfig][7] ;
  input [3:0]\slvo[11][hindex] ;
  input \slvo[10][hready] ;
  input [1:0]\slvo[10][hresp] ;
  input [31:0]\slvo[10][hrdata] ;
  input [15:0]\slvo[10][hsplit] ;
  input [31:0]\slvo[10][hirq] ;
  input [31:0]\slvo[10][hconfig][0] ;
  input [31:0]\slvo[10][hconfig][1] ;
  input [31:0]\slvo[10][hconfig][2] ;
  input [31:0]\slvo[10][hconfig][3] ;
  input [31:0]\slvo[10][hconfig][4] ;
  input [31:0]\slvo[10][hconfig][5] ;
  input [31:0]\slvo[10][hconfig][6] ;
  input [31:0]\slvo[10][hconfig][7] ;
  input [3:0]\slvo[10][hindex] ;
  input \slvo[9][hready] ;
  input [1:0]\slvo[9][hresp] ;
  input [31:0]\slvo[9][hrdata] ;
  input [15:0]\slvo[9][hsplit] ;
  input [31:0]\slvo[9][hirq] ;
  input [31:0]\slvo[9][hconfig][0] ;
  input [31:0]\slvo[9][hconfig][1] ;
  input [31:0]\slvo[9][hconfig][2] ;
  input [31:0]\slvo[9][hconfig][3] ;
  input [31:0]\slvo[9][hconfig][4] ;
  input [31:0]\slvo[9][hconfig][5] ;
  input [31:0]\slvo[9][hconfig][6] ;
  input [31:0]\slvo[9][hconfig][7] ;
  input [3:0]\slvo[9][hindex] ;
  input \slvo[8][hready] ;
  input [1:0]\slvo[8][hresp] ;
  input [31:0]\slvo[8][hrdata] ;
  input [15:0]\slvo[8][hsplit] ;
  input [31:0]\slvo[8][hirq] ;
  input [31:0]\slvo[8][hconfig][0] ;
  input [31:0]\slvo[8][hconfig][1] ;
  input [31:0]\slvo[8][hconfig][2] ;
  input [31:0]\slvo[8][hconfig][3] ;
  input [31:0]\slvo[8][hconfig][4] ;
  input [31:0]\slvo[8][hconfig][5] ;
  input [31:0]\slvo[8][hconfig][6] ;
  input [31:0]\slvo[8][hconfig][7] ;
  input [3:0]\slvo[8][hindex] ;
  input [1:0]\slvo[7][hresp] ;
  input [31:0]\slvo[7][hrdata] ;
  input [15:0]\slvo[7][hsplit] ;
  input [31:0]\slvo[7][hirq] ;
  input [31:0]\slvo[7][hconfig][0] ;
  input [31:0]\slvo[7][hconfig][1] ;
  input [31:0]\slvo[7][hconfig][2] ;
  input [31:0]\slvo[7][hconfig][3] ;
  input [31:0]\slvo[7][hconfig][4] ;
  input [31:0]\slvo[7][hconfig][5] ;
  input [31:0]\slvo[7][hconfig][6] ;
  input [31:0]\slvo[7][hconfig][7] ;
  input [3:0]\slvo[7][hindex] ;
  input \slvo[6][hready] ;
  input [1:0]\slvo[6][hresp] ;
  input [31:0]\slvo[6][hrdata] ;
  input [15:0]\slvo[6][hsplit] ;
  input [31:0]\slvo[6][hirq] ;
  input [31:0]\slvo[6][hconfig][0] ;
  input [31:0]\slvo[6][hconfig][1] ;
  input [31:0]\slvo[6][hconfig][2] ;
  input [31:0]\slvo[6][hconfig][3] ;
  input [31:0]\slvo[6][hconfig][4] ;
  input [31:0]\slvo[6][hconfig][5] ;
  input [31:0]\slvo[6][hconfig][6] ;
  input [31:0]\slvo[6][hconfig][7] ;
  input [3:0]\slvo[6][hindex] ;
  input \slvo[5][hready] ;
  input [1:0]\slvo[5][hresp] ;
  input [31:0]\slvo[5][hrdata] ;
  input [15:0]\slvo[5][hsplit] ;
  input [31:0]\slvo[5][hirq] ;
  input [31:0]\slvo[5][hconfig][0] ;
  input [31:0]\slvo[5][hconfig][1] ;
  input [31:0]\slvo[5][hconfig][2] ;
  input [31:0]\slvo[5][hconfig][3] ;
  input [31:0]\slvo[5][hconfig][4] ;
  input [31:0]\slvo[5][hconfig][5] ;
  input [31:0]\slvo[5][hconfig][6] ;
  input [31:0]\slvo[5][hconfig][7] ;
  input [3:0]\slvo[5][hindex] ;
  input \slvo[4][hready] ;
  input [1:0]\slvo[4][hresp] ;
  input [31:0]\slvo[4][hrdata] ;
  input [15:0]\slvo[4][hsplit] ;
  input [31:0]\slvo[4][hirq] ;
  input [31:0]\slvo[4][hconfig][0] ;
  input [31:0]\slvo[4][hconfig][1] ;
  input [31:0]\slvo[4][hconfig][2] ;
  input [31:0]\slvo[4][hconfig][3] ;
  input [31:0]\slvo[4][hconfig][4] ;
  input [31:0]\slvo[4][hconfig][5] ;
  input [31:0]\slvo[4][hconfig][6] ;
  input [31:0]\slvo[4][hconfig][7] ;
  input [3:0]\slvo[4][hindex] ;
  input \slvo[3][hready] ;
  input [1:0]\slvo[3][hresp] ;
  input [31:0]\slvo[3][hrdata] ;
  input [15:0]\slvo[3][hsplit] ;
  input [31:0]\slvo[3][hirq] ;
  input [31:0]\slvo[3][hconfig][0] ;
  input [31:0]\slvo[3][hconfig][1] ;
  input [31:0]\slvo[3][hconfig][2] ;
  input [31:0]\slvo[3][hconfig][3] ;
  input [31:0]\slvo[3][hconfig][4] ;
  input [31:0]\slvo[3][hconfig][5] ;
  input [31:0]\slvo[3][hconfig][6] ;
  input [31:0]\slvo[3][hconfig][7] ;
  input [3:0]\slvo[3][hindex] ;
  input \slvo[2][hready] ;
  input [1:0]\slvo[2][hresp] ;
  input [31:0]\slvo[2][hrdata] ;
  input [15:0]\slvo[2][hsplit] ;
  input [31:0]\slvo[2][hirq] ;
  input [31:0]\slvo[2][hconfig][0] ;
  input [31:0]\slvo[2][hconfig][1] ;
  input [31:0]\slvo[2][hconfig][2] ;
  input [31:0]\slvo[2][hconfig][3] ;
  input [31:0]\slvo[2][hconfig][4] ;
  input [31:0]\slvo[2][hconfig][5] ;
  input [31:0]\slvo[2][hconfig][6] ;
  input [31:0]\slvo[2][hconfig][7] ;
  input [3:0]\slvo[2][hindex] ;
  input \slvo[1][hready] ;
  input [1:0]\slvo[1][hresp] ;
  input [31:0]\slvo[1][hrdata] ;
  input [15:0]\slvo[1][hsplit] ;
  input [31:0]\slvo[1][hirq] ;
  input [31:0]\slvo[1][hconfig][0] ;
  input [31:0]\slvo[1][hconfig][1] ;
  input [31:0]\slvo[1][hconfig][2] ;
  input [31:0]\slvo[1][hconfig][3] ;
  input [31:0]\slvo[1][hconfig][4] ;
  input [31:0]\slvo[1][hconfig][5] ;
  input [31:0]\slvo[1][hconfig][6] ;
  input [31:0]\slvo[1][hconfig][7] ;
  input [3:0]\slvo[1][hindex] ;
  input \slvo[0][hready] ;
  input [1:0]\slvo[0][hresp] ;
  input [31:0]\slvo[0][hrdata] ;
  input [15:0]\slvo[0][hsplit] ;
  input [31:0]\slvo[0][hirq] ;
  input [31:0]\slvo[0][hconfig][0] ;
  input [31:0]\slvo[0][hconfig][1] ;
  input [31:0]\slvo[0][hconfig][2] ;
  input [31:0]\slvo[0][hconfig][3] ;
  input [31:0]\slvo[0][hconfig][4] ;
  input [31:0]\slvo[0][hconfig][5] ;
  input [31:0]\slvo[0][hconfig][6] ;
  input [31:0]\slvo[0][hconfig][7] ;
  input [3:0]\slvo[0][hindex] ;
  input testen;
  input testrst;
  input scanen;
  input testoen;
  input [1:0]testsig;
  input msto;
  input slvo;

  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const1>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire arb;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire arb1_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire clk;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel1166_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel1169_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel1171_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel1173_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel1192_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel2102_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel2105_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel2108_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel2119_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel2122_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel2125_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel2128_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel2139_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel2142_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel2145_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel2148_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel2159_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel2162_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel2168_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel219_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel221_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel224_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel227_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel239_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel242_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel245_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel248_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel259_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel262_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel265_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel268_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel279_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel282_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel285_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel288_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel299_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel30_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel310_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel311_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel312_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel313_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel314_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel315_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel316_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel317_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel318_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel319_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel31_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel320_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel321_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel322_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel323_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel324_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel325_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel326_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel327_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel328_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel329_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel32_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel330_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel330_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel331_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel332_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel333_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel334_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel335_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel336_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel337_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel338_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel339_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel33_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel340_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel341_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel342_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel343_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel344_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel345_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel346_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel347_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel348_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel349_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel34_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel350_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel351_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel352_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel353_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel354_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel355_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel356_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel357_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel358_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel359_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel35_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel360_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel361_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel362_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel36_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel37_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel38_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hsel39_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire msti;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:7]\^msti[hgrant] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hgrant][0]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msti[hrdata] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][0]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][0]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][0]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][10]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][10]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][10]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][11]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][11]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][11]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][12]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][12]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][12]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][13]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][13]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][13]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][14]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][14]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][14]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][15]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][15]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][15]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][16]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][16]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][16]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][17]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][17]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][17]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][18]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][18]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][18]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][19]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][19]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][19]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][1]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][1]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][1]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][20]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][20]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][20]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][21]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][21]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][21]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][22]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][22]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][22]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][23]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][23]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][23]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][24]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][24]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][24]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][25]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][25]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][25]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][26]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][26]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][26]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][27]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][27]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][27]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][28]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][28]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][28]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][29]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][29]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][29]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][2]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][2]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][2]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][30]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][30]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][30]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][31]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][31]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][31]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][3]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][3]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][3]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][4]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][4]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][4]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][5]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][5]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][5]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][6]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][6]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][6]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][7]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][7]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][7]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][8]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][8]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][8]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][9]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][9]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hrdata][9]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\msti[hresp] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hresp][0]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hresp][0]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hresp][0]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hresp][1]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msti[hresp][1]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire msto;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[0][haddr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\msto[0][hburst] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msto[0][hbusreq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[0][hconfig][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[0][hirq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msto[0][hlock] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\msto[0][hprot] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\msto[0][hsize] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\msto[0][htrans] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[0][hwdata] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msto[0][hwrite] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[1][haddr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\msto[1][hburst] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msto[1][hbusreq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[1][hconfig][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[1][hirq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msto[1][hlock] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\msto[1][hprot] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\msto[1][hsize] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\msto[1][htrans] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[1][hwdata] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msto[1][hwrite] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[2][haddr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\msto[2][hburst] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msto[2][hbusreq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[2][hconfig][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[2][hirq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msto[2][hlock] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\msto[2][hprot] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\msto[2][hsize] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\msto[2][htrans] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[2][hwdata] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msto[2][hwrite] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[3][haddr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\msto[3][hburst] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msto[3][hbusreq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[3][hconfig][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[3][hirq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msto[3][hlock] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\msto[3][hprot] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\msto[3][hsize] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\msto[3][htrans] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[3][hwdata] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msto[3][hwrite] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[4][haddr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\msto[4][hburst] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msto[4][hbusreq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[4][hconfig][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[4][hirq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msto[4][hlock] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\msto[4][hprot] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\msto[4][hsize] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\msto[4][htrans] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[4][hwdata] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msto[4][hwrite] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[5][haddr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\msto[5][hburst] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msto[5][hbusreq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[5][hconfig][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[5][hirq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msto[5][hlock] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\msto[5][hprot] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\msto[5][hsize] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\msto[5][htrans] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[5][hwdata] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msto[5][hwrite] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[6][haddr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\msto[6][hburst] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msto[6][hbusreq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[6][hconfig][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[6][hirq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msto[6][hlock] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\msto[6][hprot] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\msto[6][hsize] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\msto[6][htrans] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[6][hwdata] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msto[6][hwrite] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[7][haddr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\msto[7][hburst] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[7][hconfig][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msto[7][hlock] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\msto[7][hprot] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\msto[7][hsize] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\msto[7][htrans] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\msto[7][hwdata] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \msto[7][hwrite] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_0_in186_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_0_in5_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_11_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_14_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_179_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_185_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_1_in10_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_1_in13_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_2_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_2_in7_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_6_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rin;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rst;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire scanen;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [6:1]sel0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire slvi;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvi[haddr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][0]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][0]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][10]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][10]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][11]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][11]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][12]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][12]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][13]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][13]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][14]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][14]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][15]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][15]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][16]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][16]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][17]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][17]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][18]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][18]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][19]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][19]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][1]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][1]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][20]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][20]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][21]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][21]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][22]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][22]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][23]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][23]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][24]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][24]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][25]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][25]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][26]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][26]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][27]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][27]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][28]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][28]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][29]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][29]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][2]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][2]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][30]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][30]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][31]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][31]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][3]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][3]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][4]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][4]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][5]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][5]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][6]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][6]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][7]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][7]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][8]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][8]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][9]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[haddr][9]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\slvi[hburst] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hburst][0]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hburst][0]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hburst][1]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hburst][1]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hburst][2]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hburst][2]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvi[hirq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][0]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][0]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][10]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][10]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][11]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][11]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][12]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][12]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][13]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][13]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][14]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][14]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][15]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][15]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][16]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][16]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][17]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][17]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][18]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][18]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][19]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][19]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][1]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][1]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][20]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][20]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][21]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][21]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][22]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][22]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][23]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][23]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][24]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][24]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][25]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][25]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][26]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][26]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][27]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][27]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][28]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][28]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][29]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][29]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][2]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][2]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][30]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][30]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][31]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][31]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][3]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][3]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][4]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][4]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][5]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][5]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][6]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][6]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][7]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][7]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][8]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][8]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][9]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hirq][9]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\^slvi[hmaster] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmastlock] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [0:3]\slvi[hmbsel] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_100_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_101_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_102_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_103_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_104_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_105_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_106_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_107_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_108_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_109_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_110_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_111_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_112_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_113_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_114_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_115_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_116_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_117_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_118_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_14_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_14_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_14_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_16_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_16_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_16_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_17_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_17_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_17_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_19_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_19_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_19_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_20_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_20_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_20_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_22_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_22_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_22_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_23_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_23_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_23_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_25_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_25_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_25_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_26_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_26_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_26_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_28_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_28_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_28_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_52_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_53_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_54_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_55_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_57_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_58_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_59_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_60_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_61_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_62_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_63_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_64_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_65_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_66_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_67_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_68_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_69_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_70_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_71_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_72_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_73_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_74_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_75_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_76_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_77_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_78_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_79_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_80_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_81_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_82_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_83_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_84_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_85_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_86_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_87_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_88_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_89_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_90_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_91_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_92_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_93_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_94_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_95_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_96_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_97_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_98_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][0]_INST_0_i_99_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_100_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_101_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_102_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_103_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_104_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_105_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_106_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_107_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_108_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_109_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_110_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_111_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_112_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_113_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_114_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_115_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_116_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_12_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_12_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_12_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_14_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_14_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_14_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_15_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_15_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_15_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_17_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_17_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_17_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_18_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_18_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_18_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_20_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_20_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_20_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_21_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_21_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_21_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_23_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_23_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_23_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_24_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_24_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_24_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_26_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_26_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_26_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_52_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_53_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_54_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_55_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_57_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_58_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_59_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_60_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_61_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_62_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_63_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_64_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_65_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_66_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_67_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_68_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_69_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_70_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_71_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_72_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_73_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_74_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_75_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_76_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_77_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_78_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_79_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_80_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_81_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_82_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_83_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_84_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_85_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_86_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_87_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_88_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_89_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_90_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_91_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_92_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_93_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_94_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_95_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_96_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_97_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_98_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_99_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][1]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_26_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_26_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_26_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_28_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_28_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_28_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_29_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_29_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_29_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_31_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_31_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_31_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_32_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_32_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_34_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_34_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_34_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_52_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_53_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_54_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_55_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_57_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_58_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_59_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_60_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_61_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_62_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_63_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_64_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_65_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_66_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_67_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_68_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_69_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_6_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_6_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_6_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_70_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_71_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_72_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_73_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_74_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_75_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_76_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_77_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_78_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_79_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_80_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_81_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_82_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_83_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_84_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_85_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_86_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_87_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_88_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_89_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_8_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_8_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_90_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_91_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_92_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_93_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_94_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_95_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_96_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][2]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_12_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_12_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_12_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_9_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_9_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hmbsel][3]_INST_0_i_9_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\slvi[hprot] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hprot][0]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hprot][0]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hprot][1]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hprot][1]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hprot][2]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hprot][2]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hprot][3]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hprot][3]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hready] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hready]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hready]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hready]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [0:7]\^slvi[hsel] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_11_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_11_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_11_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_13_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_13_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_13_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_15_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_15_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_15_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_19_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_19_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_19_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_20_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_20_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_20_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_21_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_21_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_21_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_23_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_23_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_23_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_52_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_53_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_54_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_55_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_57_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_58_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_59_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_60_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_61_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_62_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_63_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_64_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_65_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_66_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_67_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_68_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_69_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_70_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_71_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_72_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_73_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_74_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_75_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_76_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_77_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_78_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_79_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_80_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_81_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_82_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_83_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_84_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_85_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_86_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_87_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_88_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_89_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_8_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_8_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_90_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_91_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_92_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][0]_INST_0_i_93_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_11_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_11_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_11_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_13_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_13_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_13_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_14_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_14_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_14_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_16_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_16_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_16_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_17_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_17_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_17_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_19_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_19_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_19_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_52_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_53_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_54_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_55_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_57_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_58_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_59_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_60_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_61_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_62_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_63_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_64_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_65_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_66_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_67_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_68_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_69_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_70_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_71_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_72_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_73_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_74_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_75_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_76_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_77_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_78_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_79_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_80_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_81_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_82_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_83_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_84_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_85_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_86_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_87_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_88_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_89_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_8_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_8_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_90_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][1]_INST_0_i_91_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_11_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_11_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_11_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_12_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_12_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_12_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_14_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_14_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_14_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_15_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_15_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_15_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_17_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_17_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_17_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_18_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_18_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_18_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_20_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_20_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_20_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_52_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_53_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_54_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_55_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_57_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_58_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_59_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_60_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_61_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_62_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_63_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_64_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_65_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_66_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_67_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_68_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_69_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_70_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_71_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_72_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_73_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_74_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_75_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_76_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_77_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_78_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_79_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_80_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_81_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_82_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_83_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_84_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_85_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_86_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_87_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_88_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_89_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_90_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_91_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_92_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_9_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_9_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][2]_INST_0_i_9_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_5_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_5_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_5_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_8_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][3]_INST_0_i_8_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_5_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_5_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_5_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][4]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][5]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][6]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_4_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_6_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_6_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_6_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsel][7]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\slvi[hsize] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsize][0]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsize][0]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsize][1]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsize][1]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsize][2]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hsize][2]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\slvi[htrans] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[htrans][0]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[htrans][0]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[htrans][1]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[htrans][1]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvi[hwdata] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][0]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][0]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][10]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][10]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][11]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][11]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][12]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][12]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][13]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][13]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][14]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][14]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][15]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][15]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][16]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][16]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][17]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][17]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][18]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][18]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][19]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][19]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][1]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][1]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][20]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][20]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][21]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][21]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][22]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][22]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][23]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][23]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][24]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][24]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][25]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][25]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][26]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][26]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][27]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][27]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][28]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][28]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][29]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][29]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][2]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][2]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][30]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][30]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][31]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][31]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][3]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][3]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][4]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][4]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][5]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][5]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][6]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][6]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][7]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][7]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][8]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][8]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][9]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwdata][9]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwrite] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwrite]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvi[hwrite]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:2]\^slvi[testin] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire slvo;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[0][hconfig][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[0][hconfig][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[0][hconfig][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[0][hconfig][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[0][hconfig][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[0][hconfig][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[0][hconfig][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[0][hconfig][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[0][hirq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[0][hrdata] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvo[0][hready] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\slvo[0][hresp] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[15][hready]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[1][hconfig][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[1][hconfig][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[1][hconfig][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[1][hconfig][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[1][hconfig][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[1][hconfig][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[1][hconfig][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[1][hconfig][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[1][hirq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[1][hrdata] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvo[1][hready] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\slvo[1][hresp] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[2][hconfig][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[2][hconfig][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[2][hconfig][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[2][hconfig][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[2][hconfig][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[2][hconfig][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[2][hconfig][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[2][hconfig][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[2][hirq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[2][hrdata] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvo[2][hready] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\slvo[2][hresp] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[3][hconfig][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[3][hconfig][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[3][hconfig][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[3][hconfig][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[3][hconfig][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[3][hconfig][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[3][hconfig][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[3][hconfig][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[3][hirq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[3][hrdata] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvo[3][hready] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\slvo[3][hresp] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[4][hconfig][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[4][hconfig][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[4][hconfig][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[4][hconfig][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[4][hconfig][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[4][hconfig][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[4][hconfig][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[4][hconfig][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[4][hirq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[4][hrdata] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvo[4][hready] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\slvo[4][hresp] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[5][hconfig][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[5][hconfig][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[5][hconfig][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[5][hconfig][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[5][hconfig][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[5][hconfig][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[5][hconfig][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[5][hconfig][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[5][hirq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[5][hrdata] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvo[5][hready] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\slvo[5][hresp] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[6][hconfig][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[6][hconfig][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[6][hconfig][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[6][hconfig][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[6][hconfig][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[6][hconfig][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[6][hconfig][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[6][hconfig][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[6][hirq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[6][hrdata] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \slvo[6][hready] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\slvo[6][hresp] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[7][hconfig][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[7][hconfig][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[7][hconfig][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[7][hconfig][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[7][hconfig][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[7][hconfig][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[7][hconfig][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[7][hconfig][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[7][hirq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\slvo[7][hrdata] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\slvo[7][hresp] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hmaster][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hmaster][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hmaster][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hmaster][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hmaster][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hmasterlock]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hmasterlock]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hmasterlock]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hmasterlock]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hmasterlock]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hmasterlock]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hmasterlockd]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][10]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][13]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][14]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][16]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][16]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][17]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][17]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][18]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][18]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][19]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][19]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][20]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][20]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][21]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][21]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][22]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][22]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][23]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][23]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][24]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][24]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][25]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][25]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][26]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][26]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][27]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][27]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][28]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][28]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][29]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][29]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][30]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][30]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatam][9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][0]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][0]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][0]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][0]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][0]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][0]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][0]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][0]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][0]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][0]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][0]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][0]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][0]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][0]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][0]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][0]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][10]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][10]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][10]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][10]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][10]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][10]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][10]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][10]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][10]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][10]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][10]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][10]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][10]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][10]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][10]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][10]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][11]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][11]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][11]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][11]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][11]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][11]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][11]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][11]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][11]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][11]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][11]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][11]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][11]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][11]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][11]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][11]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][12]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][12]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][12]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][12]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][12]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][12]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][12]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][12]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][12]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][12]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][12]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][12]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][12]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][12]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][12]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][12]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][13]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][13]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][13]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][13]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][13]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][13]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][13]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][13]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][13]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][13]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][13]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][13]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][13]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][13]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][13]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][13]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][14]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][14]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][14]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][14]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][14]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][14]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][14]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][14]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][14]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][14]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][14]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][14]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][14]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][14]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][14]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][14]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][15]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][15]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][15]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][15]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][15]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][15]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][15]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][15]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][15]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][15]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][15]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][15]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][15]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][15]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][15]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][15]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][16]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][16]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][16]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][16]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][16]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][16]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][16]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][16]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][16]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][16]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][16]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][16]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][16]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][16]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][16]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][16]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][17]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][17]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][17]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][17]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][17]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][17]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][17]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][17]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][17]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][17]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][17]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][17]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][17]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][17]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][17]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][17]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][18]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][18]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][18]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][18]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][18]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][18]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][18]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][18]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][18]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][18]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][18]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][18]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][18]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][18]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][18]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][18]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][19]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][19]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][19]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][19]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][19]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][19]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][19]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][19]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][19]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][19]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][19]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][19]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][19]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][19]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][19]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][19]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][1]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][1]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][1]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][1]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][1]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][1]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][1]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][1]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][1]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][1]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][1]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][1]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][1]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][1]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][1]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][1]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][20]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][20]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][20]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][20]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][20]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][20]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][20]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][20]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][20]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][20]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][20]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][20]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][20]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][20]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][20]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][20]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][21]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][21]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][21]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][21]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][21]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][21]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][21]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][21]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][21]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][21]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][21]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][21]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][21]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][21]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][21]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][21]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][22]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][22]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][22]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][22]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][22]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][22]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][22]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][22]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][22]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][22]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][22]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][22]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][22]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][22]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][22]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][22]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][23]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][23]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][23]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][23]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][23]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][23]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][23]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][23]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][23]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][23]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][23]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][23]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][23]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][23]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][23]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][23]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][24]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][24]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][24]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][24]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][24]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][24]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][24]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][24]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][24]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][24]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][24]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][24]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][24]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][24]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][24]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][24]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][25]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][25]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][25]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][25]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][25]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][25]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][25]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][25]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][25]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][25]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][25]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][25]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][25]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][25]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][25]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][25]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][26]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][26]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][26]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][26]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][26]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][26]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][26]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][26]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][26]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][26]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][26]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][26]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][26]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][26]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][26]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][26]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][27]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][27]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][27]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][27]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][27]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][27]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][27]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][27]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][27]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][27]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][27]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][27]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][27]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][27]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][27]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][27]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][28]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][28]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][28]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][28]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][28]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][28]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][28]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][28]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][28]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][28]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][28]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][28]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][28]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][28]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][28]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][28]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][29]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][29]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][29]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][29]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][29]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][29]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][29]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][29]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][29]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][29]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][29]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][29]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][29]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][29]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][29]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][29]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][2]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][2]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][2]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][2]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][2]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][2]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][2]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][2]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][2]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][2]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][2]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][2]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][2]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][2]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][2]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][2]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][30]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][30]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][30]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][30]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][30]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][30]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][30]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][30]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][30]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][30]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][30]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][30]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][30]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][30]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][30]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][30]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][31]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][31]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][31]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][31]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][31]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][31]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][31]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][31]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][31]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][31]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][31]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][31]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][31]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][31]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][31]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][31]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][3]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][3]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][3]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][3]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][3]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][3]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][3]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][3]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][3]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][3]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][3]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][3]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][3]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][3]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][3]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][3]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][4]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][4]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][4]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][4]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][4]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][4]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][4]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][4]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][4]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][4]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][4]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][4]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][4]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][4]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][4]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][4]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][5]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][5]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][5]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][5]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][5]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][5]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][5]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][5]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][5]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][5]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][5]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][5]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][5]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][5]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][5]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][5]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][6]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][6]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][6]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][6]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][6]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][6]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][6]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][6]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][6]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][6]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][6]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][6]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][6]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][6]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][6]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][6]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][7]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][7]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][7]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][7]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][7]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][7]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][7]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][7]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][7]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][7]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][7]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][7]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][7]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][7]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][7]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][7]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][8]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][8]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][8]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][8]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][8]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][8]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][8]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][8]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][8]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][8]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][8]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][8]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][8]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][8]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][8]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][8]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][9]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][9]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][9]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][9]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][9]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][9]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][9]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][9]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][9]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][9]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][9]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][9]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][9]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][9]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][9]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[hrdatas][9]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r[htrans][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[cfgsel_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[defslv]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[haddr][5]_rep__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[haddr][5]_rep__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[haddr][5]_rep__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[haddr][5]_rep__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[haddr][5]_rep_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[haddr][6]_rep__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[haddr][6]_rep__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[haddr][6]_rep__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[haddr][6]_rep__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[haddr][6]_rep_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[haddr][7]_rep__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[haddr][7]_rep_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[haddr_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[haddr_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[haddr_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\syncrregs.r_reg[hmasterd]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hmasterlock]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hmasterlockd]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][18]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][22]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][26]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][30]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatam][9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\syncrregs.r_reg[hrdatam]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][0]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][0]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][0]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][0]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][10]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][10]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][10]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][10]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][10]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][10]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][10]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][10]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][10]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][10]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][10]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][11]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][11]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][11]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][11]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][11]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][11]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][11]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][11]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][11]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][12]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][12]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][12]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][12]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][12]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][12]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][12]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][12]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][12]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][13]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][13]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][13]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][13]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][13]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][13]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][13]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][13]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][13]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][13]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][13]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][14]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][14]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][14]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][14]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][14]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][14]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][14]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][14]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][14]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][14]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][14]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][15]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][15]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][15]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][15]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][15]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][15]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][15]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][15]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][15]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][16]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][16]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][16]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][16]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][16]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][16]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][16]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][16]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][16]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][16]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][16]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][16]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][17]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][17]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][17]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][17]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][17]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][17]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][17]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][17]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][17]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][17]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][17]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][17]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][18]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][18]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][18]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][18]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][18]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][18]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][18]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][18]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][18]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][18]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][18]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][18]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][19]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][19]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][19]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][19]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][19]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][19]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][19]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][19]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][19]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][19]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][19]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][19]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][1]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][1]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][1]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][1]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][1]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][1]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][20]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][20]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][20]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][20]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][20]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][20]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][20]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][20]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][20]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][20]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][20]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][20]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][21]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][21]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][21]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][21]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][21]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][21]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][21]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][21]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][21]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][21]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][21]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][21]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][22]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][22]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][22]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][22]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][22]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][22]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][22]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][22]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][22]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][22]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][22]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][22]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][23]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][23]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][23]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][23]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][23]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][23]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][23]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][23]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][23]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][23]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][23]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][23]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][24]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][24]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][24]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][24]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][24]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][24]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][24]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][24]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][24]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][24]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][24]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][24]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][25]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][25]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][25]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][25]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][25]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][25]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][25]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][25]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][25]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][25]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][25]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][25]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][26]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][26]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][26]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][26]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][26]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][26]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][26]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][26]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][26]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][26]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][26]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][26]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][27]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][27]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][27]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][27]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][27]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][27]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][27]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][27]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][27]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][27]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][27]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][27]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][28]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][28]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][28]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][28]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][28]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][28]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][28]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][28]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][28]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][28]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][28]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][28]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][29]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][29]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][29]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][29]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][29]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][29]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][29]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][29]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][29]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][29]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][29]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][29]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][2]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][2]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][2]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][2]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][2]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][2]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][2]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][30]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][30]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][30]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][30]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][30]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][30]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][30]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][30]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][30]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][30]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][30]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][30]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][31]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][31]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][31]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][31]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][31]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][31]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][31]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][31]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][31]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][31]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][31]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][31]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][3]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][3]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][3]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][3]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][4]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][4]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][4]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][4]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][4]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][4]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][4]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][4]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][5]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][5]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][5]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][5]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][5]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][5]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][5]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][5]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][5]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][6]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][6]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][6]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][6]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][6]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][6]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][6]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][6]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][6]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][7]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][7]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][7]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][7]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][7]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][7]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][7]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][7]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][7]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][8]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][8]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][8]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][8]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][8]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][8]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][8]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][8]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][9]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][9]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][9]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][9]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][9]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][9]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][9]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][9]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][9]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hrdatas][9]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\syncrregs.r_reg[hrdatas]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[hready_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\syncrregs.r_reg[hslave]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \syncrregs.r_reg[htrans_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire testen;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire testoen;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire testrst;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]testsig;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire v;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:12]\v[hrdatas] ;

  assign \msti[hgrant] [0] = msti;
  assign \msti[hgrant] [1:7] = \^msti[hgrant] [1:7];
  assign \msti[hgrant] [8] = slvi;
  assign \msti[hgrant] [9] = slvi;
  assign \msti[hgrant] [10] = slvi;
  assign \msti[hgrant] [11] = slvi;
  assign \msti[hgrant] [12] = slvi;
  assign \msti[hgrant] [13] = slvi;
  assign \msti[hgrant] [14] = slvi;
  assign \msti[hgrant] [15] = slvi;
  assign \msti[hirq] [31:0] = \slvi[hirq] ;
  assign \msti[hready]  = \slvi[hready] ;
  assign \msti[scanen]  = \^slvi[testin] [2];
  assign \msti[testen]  = testen;
  assign \msti[testin] [3] = testen;
  assign \msti[testin] [2] = \^slvi[testin] [2];
  assign \msti[testin] [1:0] = testsig;
  assign \msti[testoen]  = testoen;
  assign \msti[testrst]  = testrst;
  assign \slvi[hmaster] [3] = slvi;
  assign \slvi[hmaster] [2:0] = \^slvi[hmaster] [2:0];
  assign \slvi[hsel] [0:7] = \^slvi[hsel] [0:7];
  assign \slvi[hsel] [8] = slvi;
  assign \slvi[hsel] [9] = slvi;
  assign \slvi[hsel] [10] = slvi;
  assign \slvi[hsel] [11] = slvi;
  assign \slvi[hsel] [12] = slvi;
  assign \slvi[hsel] [13] = slvi;
  assign \slvi[hsel] [14] = slvi;
  assign \slvi[hsel] [15] = slvi;
  assign \slvi[scanen]  = \^slvi[testin] [2];
  assign \slvi[testen]  = testen;
  assign \slvi[testin] [3] = testen;
  assign \slvi[testin] [2] = \^slvi[testin] [2];
  assign \slvi[testin] [1:0] = testsig;
  assign \slvi[testoen]  = testoen;
  assign \slvi[testrst]  = testrst;
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND
       (.G(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC
       (.P(\<const1>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \msti[hgrant][0]_INST_0 
       (.I0(\msti[hgrant][0]_INST_0_i_1_n_0 ),
        .I1(\msti[hgrant][0]_INST_0_i_2_n_0 ),
        .I2(\msti[hgrant][0]_INST_0_i_3_n_0 ),
        .O(msti));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBBBBBBF333BBBB)) 
    \msti[hgrant][0]_INST_0_i_1 
       (.I0(\^slvi[hmaster] [1]),
        .I1(\msti[hgrant][0]_INST_0_i_4_n_0 ),
        .I2(\msti[hgrant][0]_INST_0_i_5_n_0 ),
        .I3(\msti[hgrant][0]_INST_0_i_6_n_0 ),
        .I4(arb1_out),
        .I5(\msti[hgrant][0]_INST_0_i_8_n_0 ),
        .O(\msti[hgrant][0]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAEAFAEAEFFFFFFFF)) 
    \msti[hgrant][0]_INST_0_i_10 
       (.I0(\msti[hgrant][0]_INST_0_i_17_n_0 ),
        .I1(\msti[hgrant][0]_INST_0_i_20_n_0 ),
        .I2(\msti[hgrant][0]_INST_0_i_21_n_0 ),
        .I3(\msti[hgrant][0]_INST_0_i_22_n_0 ),
        .I4(\msti[hgrant][0]_INST_0_i_23_n_0 ),
        .I5(\msti[hgrant][0]_INST_0_i_24_n_0 ),
        .O(\msti[hgrant][0]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFBFFFFFFFFFFFF)) 
    \msti[hgrant][0]_INST_0_i_11 
       (.I0(\syncrregs.r_reg[defslv]__0 ),
        .I1(p_0_in186_in),
        .I2(\syncrregs.r_reg[cfgsel_n_0_] ),
        .I3(\msti[hresp] [0]),
        .I4(\^slvi[hmaster] [2]),
        .I5(\syncrregs.r_reg[hmasterlockd]__0 ),
        .O(\msti[hgrant][0]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFD00000000)) 
    \msti[hgrant][0]_INST_0_i_12 
       (.I0(\msti[hgrant][0]_INST_0_i_25_n_0 ),
        .I1(\msti[hgrant][0]_INST_0_i_26_n_0 ),
        .I2(\msti[hgrant][0]_INST_0_i_27_n_0 ),
        .I3(\msti[hgrant][0]_INST_0_i_22_n_0 ),
        .I4(\msti[hgrant][0]_INST_0_i_23_n_0 ),
        .I5(\msti[hgrant][0]_INST_0_i_28_n_0 ),
        .O(\msti[hgrant][0]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFEEFEFFFFFFFF)) 
    \msti[hgrant][0]_INST_0_i_13 
       (.I0(\msto[1][hbusreq] ),
        .I1(\msti[hgrant][0]_INST_0_i_23_n_0 ),
        .I2(\msto[4][hbusreq] ),
        .I3(\^slvi[hmaster] [2]),
        .I4(\msto[0][hbusreq] ),
        .I5(\msti[hgrant][0]_INST_0_i_29_n_0 ),
        .O(\msti[hgrant][0]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEF)) 
    \msti[hgrant][0]_INST_0_i_14 
       (.I0(\msto[3][hbusreq] ),
        .I1(\msto[2][hbusreq] ),
        .I2(\msto[4][hbusreq] ),
        .O(\msti[hgrant][0]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000FFCD)) 
    \msti[hgrant][0]_INST_0_i_15 
       (.I0(\msto[6][hbusreq] ),
        .I1(\msto[5][hbusreq] ),
        .I2(msto),
        .I3(\msto[4][hbusreq] ),
        .I4(\msto[2][hbusreq] ),
        .I5(\msto[3][hbusreq] ),
        .O(\msti[hgrant][0]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000FCFD)) 
    \msti[hgrant][0]_INST_0_i_16 
       (.I0(\msti[hgrant][0]_INST_0_i_26_n_0 ),
        .I1(\msti[hgrant][0]_INST_0_i_23_n_0 ),
        .I2(\msti[hgrant][0]_INST_0_i_22_n_0 ),
        .I3(\msti[hgrant][0]_INST_0_i_27_n_0 ),
        .I4(\msti[hgrant][0]_INST_0_i_21_n_0 ),
        .I5(\msti[hgrant][0]_INST_0_i_20_n_0 ),
        .O(\msti[hgrant][0]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    \msti[hgrant][0]_INST_0_i_17 
       (.I0(\msto[1][hbusreq] ),
        .I1(\^slvi[hmaster] [2]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\^slvi[hmaster] [0]),
        .O(\msti[hgrant][0]_INST_0_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1111111111111D55)) 
    \msti[hgrant][0]_INST_0_i_18 
       (.I0(\slvi[htrans] [0]),
        .I1(\slvi[htrans] [1]),
        .I2(\msti[hgrant][0]_INST_0_i_30_n_0 ),
        .I3(\slvi[hburst] [0]),
        .I4(\slvi[hburst] [1]),
        .I5(\slvi[hburst] [2]),
        .O(arb));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \msti[hgrant][0]_INST_0_i_19 
       (.I0(\msto[2][hbusreq] ),
        .I1(\msto[0][hbusreq] ),
        .I2(\msti[hgrant][0]_INST_0_i_31_n_0 ),
        .I3(\msti[hgrant][0]_INST_0_i_27_n_0 ),
        .I4(\msto[1][hbusreq] ),
        .I5(\msto[3][hbusreq] ),
        .O(\msti[hgrant][0]_INST_0_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBBBBBBF333BBBB)) 
    \msti[hgrant][0]_INST_0_i_2 
       (.I0(\^slvi[hmaster] [0]),
        .I1(\msti[hgrant][0]_INST_0_i_9_n_0 ),
        .I2(\msti[hgrant][0]_INST_0_i_10_n_0 ),
        .I3(\msti[hgrant][0]_INST_0_i_6_n_0 ),
        .I4(arb1_out),
        .I5(\msti[hgrant][0]_INST_0_i_8_n_0 ),
        .O(\msti[hgrant][0]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0222)) 
    \msti[hgrant][0]_INST_0_i_20 
       (.I0(\msto[3][hbusreq] ),
        .I1(\^slvi[hmaster] [2]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\^slvi[hmaster] [0]),
        .O(\msti[hgrant][0]_INST_0_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \msti[hgrant][0]_INST_0_i_21 
       (.I0(\msto[2][hbusreq] ),
        .I1(\^slvi[hmaster] [2]),
        .I2(\^slvi[hmaster] [1]),
        .O(\msti[hgrant][0]_INST_0_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \msti[hgrant][0]_INST_0_i_22 
       (.I0(\msto[4][hbusreq] ),
        .I1(\^slvi[hmaster] [2]),
        .O(\msti[hgrant][0]_INST_0_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h222A)) 
    \msti[hgrant][0]_INST_0_i_23 
       (.I0(\msto[5][hbusreq] ),
        .I1(\^slvi[hmaster] [2]),
        .I2(\^slvi[hmaster] [0]),
        .I3(\^slvi[hmaster] [1]),
        .O(\msti[hgrant][0]_INST_0_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5D5F5D5DFFFFFFFF)) 
    \msti[hgrant][0]_INST_0_i_24 
       (.I0(\msti[hgrant][0]_INST_0_i_32_n_0 ),
        .I1(\msto[0][hbusreq] ),
        .I2(\msti[hgrant][0]_INST_0_i_27_n_0 ),
        .I3(\msto[1][hbusreq] ),
        .I4(\msto[2][hbusreq] ),
        .I5(\msti[hgrant][0]_INST_0_i_33_n_0 ),
        .O(\msti[hgrant][0]_INST_0_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFEFFFF)) 
    \msti[hgrant][0]_INST_0_i_25 
       (.I0(\msto[3][hbusreq] ),
        .I1(\msto[1][hbusreq] ),
        .I2(\msto[0][hbusreq] ),
        .I3(\msto[2][hbusreq] ),
        .I4(\msti[hgrant][0]_INST_0_i_34_n_0 ),
        .O(\msti[hgrant][0]_INST_0_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h2A)) 
    \msti[hgrant][0]_INST_0_i_26 
       (.I0(\msto[6][hbusreq] ),
        .I1(\^slvi[hmaster] [2]),
        .I2(\^slvi[hmaster] [1]),
        .O(\msti[hgrant][0]_INST_0_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2AAA)) 
    \msti[hgrant][0]_INST_0_i_27 
       (.I0(msto),
        .I1(\^slvi[hmaster] [2]),
        .I2(\^slvi[hmaster] [0]),
        .I3(\^slvi[hmaster] [1]),
        .O(\msti[hgrant][0]_INST_0_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF000FFFFFF51)) 
    \msti[hgrant][0]_INST_0_i_28 
       (.I0(\msto[2][hbusreq] ),
        .I1(\msto[1][hbusreq] ),
        .I2(\^slvi[hmaster] [0]),
        .I3(\^slvi[hmaster] [1]),
        .I4(\^slvi[hmaster] [2]),
        .I5(\msto[3][hbusreq] ),
        .O(\msti[hgrant][0]_INST_0_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEF)) 
    \msti[hgrant][0]_INST_0_i_29 
       (.I0(\msto[3][hbusreq] ),
        .I1(\msto[2][hbusreq] ),
        .I2(\msto[5][hbusreq] ),
        .O(\msti[hgrant][0]_INST_0_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBBBBBBF333BBBB)) 
    \msti[hgrant][0]_INST_0_i_3 
       (.I0(\^slvi[hmaster] [2]),
        .I1(\msti[hgrant][0]_INST_0_i_11_n_0 ),
        .I2(\msti[hgrant][0]_INST_0_i_12_n_0 ),
        .I3(\msti[hgrant][0]_INST_0_i_6_n_0 ),
        .I4(arb1_out),
        .I5(\msti[hgrant][0]_INST_0_i_8_n_0 ),
        .O(\msti[hgrant][0]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hgrant][0]_INST_0_i_30 
       (.I0(\msti[hgrant][0]_INST_0_i_35_n_0 ),
        .I1(\msti[hgrant][0]_INST_0_i_36_n_0 ),
        .O(\msti[hgrant][0]_INST_0_i_30_n_0 ),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4400000044440404)) 
    \msti[hgrant][0]_INST_0_i_31 
       (.I0(\msti[hgrant][0]_INST_0_i_23_n_0 ),
        .I1(\msti[hgrant][0]_INST_0_i_28_n_0 ),
        .I2(\msto[4][hbusreq] ),
        .I3(\^slvi[hmaster] [1]),
        .I4(\^slvi[hmaster] [2]),
        .I5(\msto[6][hbusreq] ),
        .O(\msti[hgrant][0]_INST_0_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF000FF51)) 
    \msti[hgrant][0]_INST_0_i_32 
       (.I0(\msto[4][hbusreq] ),
        .I1(\msto[2][hbusreq] ),
        .I2(\^slvi[hmaster] [1]),
        .I3(\^slvi[hmaster] [2]),
        .I4(\msto[6][hbusreq] ),
        .O(\msti[hgrant][0]_INST_0_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h55555555FFFF55FD)) 
    \msti[hgrant][0]_INST_0_i_33 
       (.I0(\msti[hgrant][0]_INST_0_i_37_n_0 ),
        .I1(msto),
        .I2(\^slvi[hmaster] [0]),
        .I3(\msto[6][hbusreq] ),
        .I4(\msto[5][hbusreq] ),
        .I5(\msto[4][hbusreq] ),
        .O(\msti[hgrant][0]_INST_0_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \msti[hgrant][0]_INST_0_i_34 
       (.I0(\^slvi[hmaster] [2]),
        .I1(msto),
        .I2(\msto[5][hbusreq] ),
        .I3(\msto[4][hbusreq] ),
        .I4(\msto[6][hbusreq] ),
        .O(\msti[hgrant][0]_INST_0_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hgrant][0]_INST_0_i_35 
       (.I0(\msto[3][hbusreq] ),
        .I1(\msto[2][hbusreq] ),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][hbusreq] ),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][hbusreq] ),
        .O(\msti[hgrant][0]_INST_0_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hgrant][0]_INST_0_i_36 
       (.I0(msto),
        .I1(\msto[6][hbusreq] ),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][hbusreq] ),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][hbusreq] ),
        .O(\msti[hgrant][0]_INST_0_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000051111111)) 
    \msti[hgrant][0]_INST_0_i_37 
       (.I0(\msto[1][hbusreq] ),
        .I1(msto),
        .I2(\^slvi[hmaster] [2]),
        .I3(\^slvi[hmaster] [0]),
        .I4(\^slvi[hmaster] [1]),
        .I5(\msto[3][hbusreq] ),
        .O(\msti[hgrant][0]_INST_0_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFBFFFFFFFFFFFF)) 
    \msti[hgrant][0]_INST_0_i_4 
       (.I0(\syncrregs.r_reg[defslv]__0 ),
        .I1(p_0_in186_in),
        .I2(\syncrregs.r_reg[cfgsel_n_0_] ),
        .I3(\msti[hresp] [0]),
        .I4(\^slvi[hmaster] [1]),
        .I5(\syncrregs.r_reg[hmasterlockd]__0 ),
        .O(\msti[hgrant][0]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000004404FFFF)) 
    \msti[hgrant][0]_INST_0_i_5 
       (.I0(\msti[hgrant][0]_INST_0_i_13_n_0 ),
        .I1(\msti[hgrant][0]_INST_0_i_14_n_0 ),
        .I2(\msti[hgrant][0]_INST_0_i_15_n_0 ),
        .I3(\^slvi[hmaster] [1]),
        .I4(\msti[hgrant][0]_INST_0_i_16_n_0 ),
        .I5(\msti[hgrant][0]_INST_0_i_17_n_0 ),
        .O(\msti[hgrant][0]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFBFF)) 
    \msti[hgrant][0]_INST_0_i_6 
       (.I0(\syncrregs.r_reg[defslv]__0 ),
        .I1(p_0_in186_in),
        .I2(\syncrregs.r_reg[cfgsel_n_0_] ),
        .I3(\syncrregs.r_reg[hmasterlockd]__0 ),
        .I4(\msti[hresp] [0]),
        .O(\msti[hgrant][0]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \msti[hgrant][0]_INST_0_i_7 
       (.I0(arb),
        .I1(\slvi[hmastlock] ),
        .O(arb1_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \msti[hgrant][0]_INST_0_i_8 
       (.I0(\msto[6][hbusreq] ),
        .I1(\msto[4][hbusreq] ),
        .I2(\msti[hgrant][0]_INST_0_i_19_n_0 ),
        .I3(\msto[5][hbusreq] ),
        .I4(msto),
        .O(\msti[hgrant][0]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFBFFFFFFFFFFFF)) 
    \msti[hgrant][0]_INST_0_i_9 
       (.I0(\syncrregs.r_reg[defslv]__0 ),
        .I1(p_0_in186_in),
        .I2(\syncrregs.r_reg[cfgsel_n_0_] ),
        .I3(\msti[hresp] [0]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\syncrregs.r_reg[hmasterlockd]__0 ),
        .O(\msti[hgrant][0]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \msti[hgrant][1]_INST_0 
       (.I0(\msti[hgrant][0]_INST_0_i_1_n_0 ),
        .I1(\msti[hgrant][0]_INST_0_i_2_n_0 ),
        .I2(\msti[hgrant][0]_INST_0_i_3_n_0 ),
        .O(\^msti[hgrant] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \msti[hgrant][2]_INST_0 
       (.I0(\msti[hgrant][0]_INST_0_i_2_n_0 ),
        .I1(\msti[hgrant][0]_INST_0_i_1_n_0 ),
        .I2(\msti[hgrant][0]_INST_0_i_3_n_0 ),
        .O(\^msti[hgrant] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \msti[hgrant][3]_INST_0 
       (.I0(\msti[hgrant][0]_INST_0_i_1_n_0 ),
        .I1(\msti[hgrant][0]_INST_0_i_2_n_0 ),
        .I2(\msti[hgrant][0]_INST_0_i_3_n_0 ),
        .O(\^msti[hgrant] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h10)) 
    \msti[hgrant][4]_INST_0 
       (.I0(\msti[hgrant][0]_INST_0_i_1_n_0 ),
        .I1(\msti[hgrant][0]_INST_0_i_2_n_0 ),
        .I2(\msti[hgrant][0]_INST_0_i_3_n_0 ),
        .O(\^msti[hgrant] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \msti[hgrant][5]_INST_0 
       (.I0(\msti[hgrant][0]_INST_0_i_1_n_0 ),
        .I1(\msti[hgrant][0]_INST_0_i_2_n_0 ),
        .I2(\msti[hgrant][0]_INST_0_i_3_n_0 ),
        .O(\^msti[hgrant] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \msti[hgrant][6]_INST_0 
       (.I0(\msti[hgrant][0]_INST_0_i_2_n_0 ),
        .I1(\msti[hgrant][0]_INST_0_i_1_n_0 ),
        .I2(\msti[hgrant][0]_INST_0_i_3_n_0 ),
        .O(\^msti[hgrant] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \msti[hgrant][7]_INST_0 
       (.I0(\msti[hgrant][0]_INST_0_i_1_n_0 ),
        .I1(\msti[hgrant][0]_INST_0_i_2_n_0 ),
        .I2(\msti[hgrant][0]_INST_0_i_3_n_0 ),
        .O(\^msti[hgrant] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][0]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [0]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [0]),
        .I3(\msti[hrdata][0]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][0]_INST_0_i_1 
       (.I0(\msti[hrdata][0]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][0]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][0]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][0]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [0]),
        .I1(\slvo[2][hrdata] [0]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [0]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [0]),
        .O(\msti[hrdata][0]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][0]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [0]),
        .I1(\slvo[6][hrdata] [0]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [0]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [0]),
        .O(\msti[hrdata][0]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][10]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [10]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [10]),
        .I3(\msti[hrdata][10]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][10]_INST_0_i_1 
       (.I0(\msti[hrdata][10]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][10]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][10]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][10]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [10]),
        .I1(\slvo[2][hrdata] [10]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [10]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [10]),
        .O(\msti[hrdata][10]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][10]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [10]),
        .I1(\slvo[6][hrdata] [10]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [10]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [10]),
        .O(\msti[hrdata][10]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][11]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [11]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [11]),
        .I3(\msti[hrdata][11]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][11]_INST_0_i_1 
       (.I0(\msti[hrdata][11]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][11]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][11]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][11]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [11]),
        .I1(\slvo[2][hrdata] [11]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [11]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [11]),
        .O(\msti[hrdata][11]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][11]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [11]),
        .I1(\slvo[6][hrdata] [11]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [11]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [11]),
        .O(\msti[hrdata][11]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][12]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [12]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [12]),
        .I3(\msti[hrdata][12]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][12]_INST_0_i_1 
       (.I0(\msti[hrdata][12]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][12]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][12]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][12]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [12]),
        .I1(\slvo[2][hrdata] [12]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [12]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [12]),
        .O(\msti[hrdata][12]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][12]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [12]),
        .I1(\slvo[6][hrdata] [12]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [12]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [12]),
        .O(\msti[hrdata][12]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][13]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [13]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [13]),
        .I3(\msti[hrdata][13]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][13]_INST_0_i_1 
       (.I0(\msti[hrdata][13]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][13]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][13]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][13]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [13]),
        .I1(\slvo[2][hrdata] [13]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [13]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [13]),
        .O(\msti[hrdata][13]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][13]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [13]),
        .I1(\slvo[6][hrdata] [13]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [13]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [13]),
        .O(\msti[hrdata][13]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][14]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [14]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [14]),
        .I3(\msti[hrdata][14]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][14]_INST_0_i_1 
       (.I0(\msti[hrdata][14]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][14]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][14]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][14]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [14]),
        .I1(\slvo[2][hrdata] [14]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [14]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [14]),
        .O(\msti[hrdata][14]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][14]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [14]),
        .I1(\slvo[6][hrdata] [14]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [14]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [14]),
        .O(\msti[hrdata][14]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][15]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [15]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [15]),
        .I3(\msti[hrdata][15]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][15]_INST_0_i_1 
       (.I0(\msti[hrdata][15]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][15]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][15]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][15]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [15]),
        .I1(\slvo[2][hrdata] [15]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [15]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [15]),
        .O(\msti[hrdata][15]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][15]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [15]),
        .I1(\slvo[6][hrdata] [15]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [15]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [15]),
        .O(\msti[hrdata][15]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][16]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [16]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [16]),
        .I3(\msti[hrdata][16]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][16]_INST_0_i_1 
       (.I0(\msti[hrdata][16]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][16]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][16]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][16]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [16]),
        .I1(\slvo[2][hrdata] [16]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [16]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [16]),
        .O(\msti[hrdata][16]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][16]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [16]),
        .I1(\slvo[6][hrdata] [16]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [16]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [16]),
        .O(\msti[hrdata][16]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][17]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [17]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [17]),
        .I3(\msti[hrdata][17]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][17]_INST_0_i_1 
       (.I0(\msti[hrdata][17]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][17]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][17]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][17]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [17]),
        .I1(\slvo[2][hrdata] [17]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [17]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [17]),
        .O(\msti[hrdata][17]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][17]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [17]),
        .I1(\slvo[6][hrdata] [17]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [17]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [17]),
        .O(\msti[hrdata][17]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][18]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [18]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [18]),
        .I3(\msti[hrdata][18]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][18]_INST_0_i_1 
       (.I0(\msti[hrdata][18]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][18]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][18]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][18]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [18]),
        .I1(\slvo[2][hrdata] [18]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [18]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [18]),
        .O(\msti[hrdata][18]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][18]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [18]),
        .I1(\slvo[6][hrdata] [18]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [18]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [18]),
        .O(\msti[hrdata][18]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][19]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [19]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [19]),
        .I3(\msti[hrdata][19]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][19]_INST_0_i_1 
       (.I0(\msti[hrdata][19]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][19]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][19]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][19]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [19]),
        .I1(\slvo[2][hrdata] [19]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [19]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [19]),
        .O(\msti[hrdata][19]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][19]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [19]),
        .I1(\slvo[6][hrdata] [19]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [19]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [19]),
        .O(\msti[hrdata][19]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][1]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [1]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [1]),
        .I3(\msti[hrdata][1]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][1]_INST_0_i_1 
       (.I0(\msti[hrdata][1]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][1]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][1]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][1]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [1]),
        .I1(\slvo[2][hrdata] [1]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [1]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [1]),
        .O(\msti[hrdata][1]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][1]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [1]),
        .I1(\slvo[6][hrdata] [1]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [1]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [1]),
        .O(\msti[hrdata][1]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][20]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [20]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [20]),
        .I3(\msti[hrdata][20]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][20]_INST_0_i_1 
       (.I0(\msti[hrdata][20]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][20]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][20]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][20]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [20]),
        .I1(\slvo[2][hrdata] [20]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [20]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [20]),
        .O(\msti[hrdata][20]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][20]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [20]),
        .I1(\slvo[6][hrdata] [20]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [20]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [20]),
        .O(\msti[hrdata][20]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][21]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [21]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [21]),
        .I3(\msti[hrdata][21]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][21]_INST_0_i_1 
       (.I0(\msti[hrdata][21]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][21]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][21]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F))
    \msti[hrdata][21]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [21]),
        .I1(\slvo[2][hrdata] [21]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [21]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [21]),
        .O(\msti[hrdata][21]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][21]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [21]),
        .I1(\slvo[6][hrdata] [21]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [21]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [21]),
        .O(\msti[hrdata][21]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][22]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [22]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [22]),
        .I3(\msti[hrdata][22]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][22]_INST_0_i_1 
       (.I0(\msti[hrdata][22]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][22]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][22]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][22]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [22]),
        .I1(\slvo[2][hrdata] [22]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [22]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [22]),
        .O(\msti[hrdata][22]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][22]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [22]),
        .I1(\slvo[6][hrdata] [22]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [22]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [22]),
        .O(\msti[hrdata][22]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][23]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [23]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [23]),
        .I3(\msti[hrdata][23]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][23]_INST_0_i_1 
       (.I0(\msti[hrdata][23]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][23]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][23]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][23]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [23]),
        .I1(\slvo[2][hrdata] [23]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [23]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [23]),
        .O(\msti[hrdata][23]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][23]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [23]),
        .I1(\slvo[6][hrdata] [23]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [23]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [23]),
        .O(\msti[hrdata][23]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][24]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [24]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [24]),
        .I3(\msti[hrdata][24]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][24]_INST_0_i_1 
       (.I0(\msti[hrdata][24]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][24]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][24]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][24]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [24]),
        .I1(\slvo[2][hrdata] [24]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [24]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [24]),
        .O(\msti[hrdata][24]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][24]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [24]),
        .I1(\slvo[6][hrdata] [24]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [24]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [24]),
        .O(\msti[hrdata][24]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][25]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [25]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [25]),
        .I3(\msti[hrdata][25]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][25]_INST_0_i_1 
       (.I0(\msti[hrdata][25]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][25]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][25]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][25]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [25]),
        .I1(\slvo[2][hrdata] [25]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [25]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [25]),
        .O(\msti[hrdata][25]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][25]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [25]),
        .I1(\slvo[6][hrdata] [25]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [25]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [25]),
        .O(\msti[hrdata][25]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][26]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [26]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [26]),
        .I3(\msti[hrdata][26]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][26]_INST_0_i_1 
       (.I0(\msti[hrdata][26]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][26]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][26]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][26]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [26]),
        .I1(\slvo[2][hrdata] [26]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [26]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [26]),
        .O(\msti[hrdata][26]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][26]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [26]),
        .I1(\slvo[6][hrdata] [26]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [26]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [26]),
        .O(\msti[hrdata][26]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][27]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [27]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [27]),
        .I3(\msti[hrdata][27]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][27]_INST_0_i_1 
       (.I0(\msti[hrdata][27]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][27]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][27]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][27]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [27]),
        .I1(\slvo[2][hrdata] [27]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [27]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [27]),
        .O(\msti[hrdata][27]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][27]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [27]),
        .I1(\slvo[6][hrdata] [27]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [27]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [27]),
        .O(\msti[hrdata][27]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][28]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [28]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [28]),
        .I3(\msti[hrdata][28]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][28]_INST_0_i_1 
       (.I0(\msti[hrdata][28]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][28]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][28]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][28]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [28]),
        .I1(\slvo[2][hrdata] [28]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [28]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [28]),
        .O(\msti[hrdata][28]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][28]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [28]),
        .I1(\slvo[6][hrdata] [28]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [28]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [28]),
        .O(\msti[hrdata][28]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][29]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [29]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [29]),
        .I3(\msti[hrdata][29]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][29]_INST_0_i_1 
       (.I0(\msti[hrdata][29]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][29]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][29]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][29]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [29]),
        .I1(\slvo[2][hrdata] [29]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [29]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [29]),
        .O(\msti[hrdata][29]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][29]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [29]),
        .I1(\slvo[6][hrdata] [29]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [29]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [29]),
        .O(\msti[hrdata][29]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][2]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [2]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [2]),
        .I3(\msti[hrdata][2]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][2]_INST_0_i_1 
       (.I0(\msti[hrdata][2]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][2]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][2]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][2]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [2]),
        .I1(\slvo[2][hrdata] [2]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [2]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [2]),
        .O(\msti[hrdata][2]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][2]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [2]),
        .I1(\slvo[6][hrdata] [2]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [2]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [2]),
        .O(\msti[hrdata][2]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][30]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [30]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [30]),
        .I3(\msti[hrdata][30]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][30]_INST_0_i_1 
       (.I0(\msti[hrdata][30]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][30]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][30]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][30]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [30]),
        .I1(\slvo[2][hrdata] [30]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [30]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [30]),
        .O(\msti[hrdata][30]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][30]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [30]),
        .I1(\slvo[6][hrdata] [30]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [30]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [30]),
        .O(\msti[hrdata][30]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][31]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [31]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [31]),
        .I3(\msti[hrdata][31]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][31]_INST_0_i_1 
       (.I0(\msti[hrdata][31]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][31]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][31]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][31]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [31]),
        .I1(\slvo[2][hrdata] [31]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [31]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [31]),
        .O(\msti[hrdata][31]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][31]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [31]),
        .I1(\slvo[6][hrdata] [31]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [31]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [31]),
        .O(\msti[hrdata][31]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][3]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [3]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [3]),
        .I3(\msti[hrdata][3]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][3]_INST_0_i_1 
       (.I0(\msti[hrdata][3]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][3]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][3]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][3]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [3]),
        .I1(\slvo[2][hrdata] [3]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [3]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [3]),
        .O(\msti[hrdata][3]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][3]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [3]),
        .I1(\slvo[6][hrdata] [3]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [3]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [3]),
        .O(\msti[hrdata][3]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][4]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [4]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [4]),
        .I3(\msti[hrdata][4]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][4]_INST_0_i_1 
       (.I0(\msti[hrdata][4]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][4]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][4]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][4]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [4]),
        .I1(\slvo[2][hrdata] [4]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [4]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [4]),
        .O(\msti[hrdata][4]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][4]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [4]),
        .I1(\slvo[6][hrdata] [4]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [4]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [4]),
        .O(\msti[hrdata][4]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][5]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [5]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [5]),
        .I3(\msti[hrdata][5]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][5]_INST_0_i_1 
       (.I0(\msti[hrdata][5]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][5]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][5]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][5]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [5]),
        .I1(\slvo[2][hrdata] [5]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [5]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [5]),
        .O(\msti[hrdata][5]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][5]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [5]),
        .I1(\slvo[6][hrdata] [5]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [5]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [5]),
        .O(\msti[hrdata][5]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][6]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [6]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [6]),
        .I3(\msti[hrdata][6]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][6]_INST_0_i_1 
       (.I0(\msti[hrdata][6]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][6]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][6]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][6]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [6]),
        .I1(\slvo[2][hrdata] [6]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [6]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [6]),
        .O(\msti[hrdata][6]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][6]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [6]),
        .I1(\slvo[6][hrdata] [6]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [6]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [6]),
        .O(\msti[hrdata][6]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][7]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [7]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [7]),
        .I3(\msti[hrdata][7]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][7]_INST_0_i_1 
       (.I0(\msti[hrdata][7]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][7]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][7]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][7]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [7]),
        .I1(\slvo[2][hrdata] [7]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [7]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [7]),
        .O(\msti[hrdata][7]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][7]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [7]),
        .I1(\slvo[6][hrdata] [7]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [7]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [7]),
        .O(\msti[hrdata][7]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][8]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [8]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [8]),
        .I3(\msti[hrdata][8]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][8]_INST_0_i_1 
       (.I0(\msti[hrdata][8]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][8]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][8]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][8]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [8]),
        .I1(\slvo[2][hrdata] [8]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [8]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [8]),
        .O(\msti[hrdata][8]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][8]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [8]),
        .I1(\slvo[6][hrdata] [8]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [8]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [8]),
        .O(\msti[hrdata][8]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \msti[hrdata][9]_INST_0 
       (.I0(\syncrregs.r_reg[hrdatas]__0 [9]),
        .I1(\syncrregs.r_reg ),
        .I2(\syncrregs.r_reg[hrdatam]__0 [9]),
        .I3(\msti[hrdata][9]_INST_0_i_1_n_0 ),
        .I4(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hrdata] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hrdata][9]_INST_0_i_1 
       (.I0(\msti[hrdata][9]_INST_0_i_2_n_0 ),
        .I1(\msti[hrdata][9]_INST_0_i_3_n_0 ),
        .O(\msti[hrdata][9]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][9]_INST_0_i_2 
       (.I0(\slvo[3][hrdata] [9]),
        .I1(\slvo[2][hrdata] [9]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hrdata] [9]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hrdata] [9]),
        .O(\msti[hrdata][9]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hrdata][9]_INST_0_i_3 
       (.I0(\slvo[7][hrdata] [9]),
        .I1(\slvo[6][hrdata] [9]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hrdata] [9]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hrdata] [9]),
        .O(\msti[hrdata][9]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00E4)) 
    \msti[hresp][0]_INST_0 
       (.I0(\syncrregs.r_reg[defslv]__0 ),
        .I1(\msti[hresp][0]_INST_0_i_1_n_0 ),
        .I2(\syncrregs.r_reg[htrans_n_0_][1] ),
        .I3(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hresp] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hresp][0]_INST_0_i_1 
       (.I0(\msti[hresp][0]_INST_0_i_2_n_0 ),
        .I1(\msti[hresp][0]_INST_0_i_3_n_0 ),
        .O(\msti[hresp][0]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hresp][0]_INST_0_i_2 
       (.I0(\slvo[3][hresp] [0]),
        .I1(\slvo[2][hresp] [0]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hresp] [0]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hresp] [0]),
        .O(\msti[hresp][0]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hresp][0]_INST_0_i_3 
       (.I0(\slvo[7][hresp] [0]),
        .I1(\slvo[6][hresp] [0]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hresp] [0]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hresp] [0]),
        .O(\msti[hresp][0]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \msti[hresp][1]_INST_0 
       (.I0(\syncrregs.r_reg[defslv]__0 ),
        .I1(p_0_in186_in),
        .I2(\syncrregs.r_reg[cfgsel_n_0_] ),
        .O(\msti[hresp] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \msti[hresp][1]_INST_0_i_1 
       (.I0(\msti[hresp][1]_INST_0_i_2_n_0 ),
        .I1(\msti[hresp][1]_INST_0_i_3_n_0 ),
        .O(p_0_in186_in),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hresp][1]_INST_0_i_2 
       (.I0(\slvo[3][hresp] [1]),
        .I1(\slvo[2][hresp] [1]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hresp] [1]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hresp] [1]),
        .O(\msti[hresp][1]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \msti[hresp][1]_INST_0_i_3 
       (.I0(\slvo[7][hresp] [1]),
        .I1(\slvo[6][hresp] [1]),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hresp] [1]),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hresp] [1]),
        .O(\msti[hresp][1]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][0]_INST_0 
       (.I0(\slvi[haddr][0]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][0]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [0]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][0]_INST_0_i_1 
       (.I0(\msto[3][haddr] [0]),
        .I1(\msto[2][haddr] [0]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [0]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [0]),
        .O(\slvi[haddr][0]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][0]_INST_0_i_2 
       (.I0(\msto[7][haddr] [0]),
        .I1(\msto[6][haddr] [0]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [0]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [0]),
        .O(\slvi[haddr][0]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][10]_INST_0 
       (.I0(\slvi[haddr][10]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][10]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [10]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][10]_INST_0_i_1 
       (.I0(\msto[3][haddr] [10]),
        .I1(\msto[2][haddr] [10]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [10]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [10]),
        .O(\slvi[haddr][10]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][10]_INST_0_i_2 
       (.I0(\msto[7][haddr] [10]),
        .I1(\msto[6][haddr] [10]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [10]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [10]),
        .O(\slvi[haddr][10]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][11]_INST_0 
       (.I0(\slvi[haddr][11]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][11]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [11]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][11]_INST_0_i_1 
       (.I0(\msto[3][haddr] [11]),
        .I1(\msto[2][haddr] [11]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [11]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [11]),
        .O(\slvi[haddr][11]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][11]_INST_0_i_2 
       (.I0(\msto[7][haddr] [11]),
        .I1(\msto[6][haddr] [11]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [11]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [11]),
        .O(\slvi[haddr][11]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][12]_INST_0 
       (.I0(\slvi[haddr][12]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][12]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [12]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][12]_INST_0_i_1 
       (.I0(\msto[3][haddr] [12]),
        .I1(\msto[2][haddr] [12]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [12]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [12]),
        .O(\slvi[haddr][12]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][12]_INST_0_i_2 
       (.I0(\msto[7][haddr] [12]),
        .I1(\msto[6][haddr] [12]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [12]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [12]),
        .O(\slvi[haddr][12]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][13]_INST_0 
       (.I0(\slvi[haddr][13]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][13]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [13]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][13]_INST_0_i_1 
       (.I0(\msto[3][haddr] [13]),
        .I1(\msto[2][haddr] [13]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [13]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [13]),
        .O(\slvi[haddr][13]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][13]_INST_0_i_2 
       (.I0(\msto[7][haddr] [13]),
        .I1(\msto[6][haddr] [13]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [13]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [13]),
        .O(\slvi[haddr][13]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][14]_INST_0 
       (.I0(\slvi[haddr][14]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][14]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [14]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][14]_INST_0_i_1 
       (.I0(\msto[3][haddr] [14]),
        .I1(\msto[2][haddr] [14]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [14]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [14]),
        .O(\slvi[haddr][14]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][14]_INST_0_i_2 
       (.I0(\msto[7][haddr] [14]),
        .I1(\msto[6][haddr] [14]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [14]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [14]),
        .O(\slvi[haddr][14]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][15]_INST_0 
       (.I0(\slvi[haddr][15]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][15]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [15]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][15]_INST_0_i_1 
       (.I0(\msto[3][haddr] [15]),
        .I1(\msto[2][haddr] [15]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [15]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [15]),
        .O(\slvi[haddr][15]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][15]_INST_0_i_2 
       (.I0(\msto[7][haddr] [15]),
        .I1(\msto[6][haddr] [15]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [15]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [15]),
        .O(\slvi[haddr][15]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][16]_INST_0 
       (.I0(\slvi[haddr][16]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][16]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [16]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][16]_INST_0_i_1 
       (.I0(\msto[3][haddr] [16]),
        .I1(\msto[2][haddr] [16]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [16]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [16]),
        .O(\slvi[haddr][16]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][16]_INST_0_i_2 
       (.I0(\msto[7][haddr] [16]),
        .I1(\msto[6][haddr] [16]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [16]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [16]),
        .O(\slvi[haddr][16]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][17]_INST_0 
       (.I0(\slvi[haddr][17]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][17]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [17]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][17]_INST_0_i_1 
       (.I0(\msto[3][haddr] [17]),
        .I1(\msto[2][haddr] [17]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [17]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [17]),
        .O(\slvi[haddr][17]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][17]_INST_0_i_2 
       (.I0(\msto[7][haddr] [17]),
        .I1(\msto[6][haddr] [17]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [17]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [17]),
        .O(\slvi[haddr][17]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][18]_INST_0 
       (.I0(\slvi[haddr][18]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][18]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [18]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][18]_INST_0_i_1 
       (.I0(\msto[3][haddr] [18]),
        .I1(\msto[2][haddr] [18]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [18]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [18]),
        .O(\slvi[haddr][18]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][18]_INST_0_i_2 
       (.I0(\msto[7][haddr] [18]),
        .I1(\msto[6][haddr] [18]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [18]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [18]),
        .O(\slvi[haddr][18]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][19]_INST_0 
       (.I0(\slvi[haddr][19]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][19]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [19]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][19]_INST_0_i_1 
       (.I0(\msto[3][haddr] [19]),
        .I1(\msto[2][haddr] [19]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [19]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [19]),
        .O(\slvi[haddr][19]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][19]_INST_0_i_2 
       (.I0(\msto[7][haddr] [19]),
        .I1(\msto[6][haddr] [19]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [19]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [19]),
        .O(\slvi[haddr][19]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][1]_INST_0 
       (.I0(\slvi[haddr][1]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][1]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [1]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][1]_INST_0_i_1 
       (.I0(\msto[3][haddr] [1]),
        .I1(\msto[2][haddr] [1]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [1]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [1]),
        .O(\slvi[haddr][1]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][1]_INST_0_i_2 
       (.I0(\msto[7][haddr] [1]),
        .I1(\msto[6][haddr] [1]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [1]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [1]),
        .O(\slvi[haddr][1]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][20]_INST_0 
       (.I0(\slvi[haddr][20]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][20]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [20]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][20]_INST_0_i_1 
       (.I0(\msto[3][haddr] [20]),
        .I1(\msto[2][haddr] [20]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [20]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [20]),
        .O(\slvi[haddr][20]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][20]_INST_0_i_2 
       (.I0(\msto[7][haddr] [20]),
        .I1(\msto[6][haddr] [20]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [20]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [20]),
        .O(\slvi[haddr][20]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][21]_INST_0 
       (.I0(\slvi[haddr][21]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][21]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [21]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][21]_INST_0_i_1 
       (.I0(\msto[3][haddr] [21]),
        .I1(\msto[2][haddr] [21]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [21]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [21]),
        .O(\slvi[haddr][21]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][21]_INST_0_i_2 
       (.I0(\msto[7][haddr] [21]),
        .I1(\msto[6][haddr] [21]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [21]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [21]),
        .O(\slvi[haddr][21]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][22]_INST_0 
       (.I0(\slvi[haddr][22]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][22]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [22]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][22]_INST_0_i_1 
       (.I0(\msto[3][haddr] [22]),
        .I1(\msto[2][haddr] [22]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [22]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [22]),
        .O(\slvi[haddr][22]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][22]_INST_0_i_2 
       (.I0(\msto[7][haddr] [22]),
        .I1(\msto[6][haddr] [22]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [22]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [22]),
        .O(\slvi[haddr][22]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][23]_INST_0 
       (.I0(\slvi[haddr][23]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][23]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [23]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][23]_INST_0_i_1 
       (.I0(\msto[3][haddr] [23]),
        .I1(\msto[2][haddr] [23]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [23]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [23]),
        .O(\slvi[haddr][23]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][23]_INST_0_i_2 
       (.I0(\msto[7][haddr] [23]),
        .I1(\msto[6][haddr] [23]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [23]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [23]),
        .O(\slvi[haddr][23]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][24]_INST_0 
       (.I0(\slvi[haddr][24]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][24]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [24]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][24]_INST_0_i_1 
       (.I0(\msto[3][haddr] [24]),
        .I1(\msto[2][haddr] [24]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [24]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [24]),
        .O(\slvi[haddr][24]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][24]_INST_0_i_2 
       (.I0(\msto[7][haddr] [24]),
        .I1(\msto[6][haddr] [24]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [24]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [24]),
        .O(\slvi[haddr][24]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][25]_INST_0 
       (.I0(\slvi[haddr][25]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][25]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [25]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][25]_INST_0_i_1 
       (.I0(\msto[3][haddr] [25]),
        .I1(\msto[2][haddr] [25]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [25]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [25]),
        .O(\slvi[haddr][25]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][25]_INST_0_i_2 
       (.I0(\msto[7][haddr] [25]),
        .I1(\msto[6][haddr] [25]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [25]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [25]),
        .O(\slvi[haddr][25]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][26]_INST_0 
       (.I0(\slvi[haddr][26]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][26]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [26]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][26]_INST_0_i_1 
       (.I0(\msto[3][haddr] [26]),
        .I1(\msto[2][haddr] [26]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [26]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [26]),
        .O(\slvi[haddr][26]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][26]_INST_0_i_2 
       (.I0(\msto[7][haddr] [26]),
        .I1(\msto[6][haddr] [26]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [26]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [26]),
        .O(\slvi[haddr][26]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][27]_INST_0 
       (.I0(\slvi[haddr][27]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][27]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [27]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][27]_INST_0_i_1 
       (.I0(\msto[3][haddr] [27]),
        .I1(\msto[2][haddr] [27]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [27]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [27]),
        .O(\slvi[haddr][27]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][27]_INST_0_i_2 
       (.I0(\msto[7][haddr] [27]),
        .I1(\msto[6][haddr] [27]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [27]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [27]),
        .O(\slvi[haddr][27]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][28]_INST_0 
       (.I0(\slvi[haddr][28]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][28]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [28]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][28]_INST_0_i_1 
       (.I0(\msto[3][haddr] [28]),
        .I1(\msto[2][haddr] [28]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [28]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [28]),
        .O(\slvi[haddr][28]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][28]_INST_0_i_2 
       (.I0(\msto[7][haddr] [28]),
        .I1(\msto[6][haddr] [28]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [28]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [28]),
        .O(\slvi[haddr][28]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][29]_INST_0 
       (.I0(\slvi[haddr][29]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][29]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [29]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][29]_INST_0_i_1 
       (.I0(\msto[3][haddr] [29]),
        .I1(\msto[2][haddr] [29]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [29]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [29]),
        .O(\slvi[haddr][29]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][29]_INST_0_i_2 
       (.I0(\msto[7][haddr] [29]),
        .I1(\msto[6][haddr] [29]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [29]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [29]),
        .O(\slvi[haddr][29]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][2]_INST_0 
       (.I0(\slvi[haddr][2]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][2]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [2]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][2]_INST_0_i_1 
       (.I0(\msto[3][haddr] [2]),
        .I1(\msto[2][haddr] [2]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [2]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [2]),
        .O(\slvi[haddr][2]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][2]_INST_0_i_2 
       (.I0(\msto[7][haddr] [2]),
        .I1(\msto[6][haddr] [2]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [2]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [2]),
        .O(\slvi[haddr][2]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][30]_INST_0 
       (.I0(\slvi[haddr][30]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][30]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [30]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][30]_INST_0_i_1 
       (.I0(\msto[3][haddr] [30]),
        .I1(\msto[2][haddr] [30]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [30]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [30]),
        .O(\slvi[haddr][30]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][30]_INST_0_i_2 
       (.I0(\msto[7][haddr] [30]),
        .I1(\msto[6][haddr] [30]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [30]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [30]),
        .O(\slvi[haddr][30]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][31]_INST_0 
       (.I0(\slvi[haddr][31]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][31]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [31]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][31]_INST_0_i_1 
       (.I0(\msto[3][haddr] [31]),
        .I1(\msto[2][haddr] [31]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [31]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [31]),
        .O(\slvi[haddr][31]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][31]_INST_0_i_2 
       (.I0(\msto[7][haddr] [31]),
        .I1(\msto[6][haddr] [31]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [31]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [31]),
        .O(\slvi[haddr][31]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][3]_INST_0 
       (.I0(\slvi[haddr][3]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][3]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [3]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][3]_INST_0_i_1 
       (.I0(\msto[3][haddr] [3]),
        .I1(\msto[2][haddr] [3]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [3]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [3]),
        .O(\slvi[haddr][3]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][3]_INST_0_i_2 
       (.I0(\msto[7][haddr] [3]),
        .I1(\msto[6][haddr] [3]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [3]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [3]),
        .O(\slvi[haddr][3]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][4]_INST_0 
       (.I0(\slvi[haddr][4]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][4]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [4]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][4]_INST_0_i_1 
       (.I0(\msto[3][haddr] [4]),
        .I1(\msto[2][haddr] [4]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [4]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [4]),
        .O(\slvi[haddr][4]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][4]_INST_0_i_2 
       (.I0(\msto[7][haddr] [4]),
        .I1(\msto[6][haddr] [4]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [4]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [4]),
        .O(\slvi[haddr][4]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][5]_INST_0 
       (.I0(\slvi[haddr][5]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][5]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [5]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][5]_INST_0_i_1 
       (.I0(\msto[3][haddr] [5]),
        .I1(\msto[2][haddr] [5]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [5]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [5]),
        .O(\slvi[haddr][5]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][5]_INST_0_i_2 
       (.I0(\msto[7][haddr] [5]),
        .I1(\msto[6][haddr] [5]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [5]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [5]),
        .O(\slvi[haddr][5]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][6]_INST_0 
       (.I0(\slvi[haddr][6]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][6]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [6]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][6]_INST_0_i_1 
       (.I0(\msto[3][haddr] [6]),
        .I1(\msto[2][haddr] [6]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [6]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [6]),
        .O(\slvi[haddr][6]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][6]_INST_0_i_2 
       (.I0(\msto[7][haddr] [6]),
        .I1(\msto[6][haddr] [6]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [6]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [6]),
        .O(\slvi[haddr][6]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][7]_INST_0 
       (.I0(\slvi[haddr][7]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][7]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [7]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][7]_INST_0_i_1 
       (.I0(\msto[3][haddr] [7]),
        .I1(\msto[2][haddr] [7]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [7]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [7]),
        .O(\slvi[haddr][7]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][7]_INST_0_i_2 
       (.I0(\msto[7][haddr] [7]),
        .I1(\msto[6][haddr] [7]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [7]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [7]),
        .O(\slvi[haddr][7]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][8]_INST_0 
       (.I0(\slvi[haddr][8]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][8]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [8]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][8]_INST_0_i_1 
       (.I0(\msto[3][haddr] [8]),
        .I1(\msto[2][haddr] [8]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [8]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [8]),
        .O(\slvi[haddr][8]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][8]_INST_0_i_2 
       (.I0(\msto[7][haddr] [8]),
        .I1(\msto[6][haddr] [8]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [8]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [8]),
        .O(\slvi[haddr][8]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[haddr][9]_INST_0 
       (.I0(\slvi[haddr][9]_INST_0_i_1_n_0 ),
        .I1(\slvi[haddr][9]_INST_0_i_2_n_0 ),
        .O(\slvi[haddr] [9]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][9]_INST_0_i_1 
       (.I0(\msto[3][haddr] [9]),
        .I1(\msto[2][haddr] [9]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][haddr] [9]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][haddr] [9]),
        .O(\slvi[haddr][9]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[haddr][9]_INST_0_i_2 
       (.I0(\msto[7][haddr] [9]),
        .I1(\msto[6][haddr] [9]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][haddr] [9]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][haddr] [9]),
        .O(\slvi[haddr][9]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hburst][0]_INST_0 
       (.I0(\slvi[hburst][0]_INST_0_i_1_n_0 ),
        .I1(\slvi[hburst][0]_INST_0_i_2_n_0 ),
        .O(\slvi[hburst] [0]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hburst][0]_INST_0_i_1 
       (.I0(\msto[3][hburst] [0]),
        .I1(\msto[2][hburst] [0]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][hburst] [0]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][hburst] [0]),
        .O(\slvi[hburst][0]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hburst][0]_INST_0_i_2 
       (.I0(\msto[7][hburst] [0]),
        .I1(\msto[6][hburst] [0]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][hburst] [0]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][hburst] [0]),
        .O(\slvi[hburst][0]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hburst][1]_INST_0 
       (.I0(\slvi[hburst][1]_INST_0_i_1_n_0 ),
        .I1(\slvi[hburst][1]_INST_0_i_2_n_0 ),
        .O(\slvi[hburst] [1]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hburst][1]_INST_0_i_1 
       (.I0(\msto[3][hburst] [1]),
        .I1(\msto[2][hburst] [1]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][hburst] [1]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][hburst] [1]),
        .O(\slvi[hburst][1]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hburst][1]_INST_0_i_2 
       (.I0(\msto[7][hburst] [1]),
        .I1(\msto[6][hburst] [1]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][hburst] [1]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][hburst] [1]),
        .O(\slvi[hburst][1]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hburst][2]_INST_0 
       (.I0(\slvi[hburst][2]_INST_0_i_1_n_0 ),
        .I1(\slvi[hburst][2]_INST_0_i_2_n_0 ),
        .O(\slvi[hburst] [2]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hburst][2]_INST_0_i_1 
       (.I0(\msto[3][hburst] [2]),
        .I1(\msto[2][hburst] [2]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][hburst] [2]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][hburst] [2]),
        .O(\slvi[hburst][2]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hburst][2]_INST_0_i_2 
       (.I0(\msto[7][hburst] [2]),
        .I1(\msto[6][hburst] [2]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][hburst] [2]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][hburst] [2]),
        .O(\slvi[hburst][2]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][0]_INST_0 
       (.I0(\slvi[hirq][0]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][0]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [0]),
        .I3(\slvo[1][hirq] [0]),
        .I4(\slvo[3][hirq] [0]),
        .O(\slvi[hirq] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][0]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [0]),
        .I1(\msto[6][hirq] [0]),
        .I2(\msto[4][hirq] [0]),
        .I3(\msto[5][hirq] [0]),
        .I4(\msto[3][hirq] [0]),
        .I5(\msto[2][hirq] [0]),
        .O(\slvi[hirq][0]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][0]_INST_0_i_2 
       (.I0(\msto[0][hirq] [0]),
        .I1(\msto[1][hirq] [0]),
        .I2(\slvo[6][hirq] [0]),
        .I3(\slvo[7][hirq] [0]),
        .I4(\slvo[5][hirq] [0]),
        .I5(\slvo[4][hirq] [0]),
        .O(\slvi[hirq][0]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][10]_INST_0 
       (.I0(\slvi[hirq][10]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][10]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [10]),
        .I3(\slvo[1][hirq] [10]),
        .I4(\slvo[3][hirq] [10]),
        .O(\slvi[hirq] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][10]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [10]),
        .I1(\msto[6][hirq] [10]),
        .I2(\msto[4][hirq] [10]),
        .I3(\msto[5][hirq] [10]),
        .I4(\msto[3][hirq] [10]),
        .I5(\msto[2][hirq] [10]),
        .O(\slvi[hirq][10]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][10]_INST_0_i_2 
       (.I0(\msto[0][hirq] [10]),
        .I1(\msto[1][hirq] [10]),
        .I2(\slvo[6][hirq] [10]),
        .I3(\slvo[7][hirq] [10]),
        .I4(\slvo[5][hirq] [10]),
        .I5(\slvo[4][hirq] [10]),
        .O(\slvi[hirq][10]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][11]_INST_0 
       (.I0(\slvi[hirq][11]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][11]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [11]),
        .I3(\slvo[1][hirq] [11]),
        .I4(\slvo[3][hirq] [11]),
        .O(\slvi[hirq] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][11]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [11]),
        .I1(\msto[6][hirq] [11]),
        .I2(\msto[4][hirq] [11]),
        .I3(\msto[5][hirq] [11]),
        .I4(\msto[3][hirq] [11]),
        .I5(\msto[2][hirq] [11]),
        .O(\slvi[hirq][11]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][11]_INST_0_i_2 
       (.I0(\msto[0][hirq] [11]),
        .I1(\msto[1][hirq] [11]),
        .I2(\slvo[6][hirq] [11]),
        .I3(\slvo[7][hirq] [11]),
        .I4(\slvo[5][hirq] [11]),
        .I5(\slvo[4][hirq] [11]),
        .O(\slvi[hirq][11]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][12]_INST_0 
       (.I0(\slvi[hirq][12]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][12]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [12]),
        .I3(\slvo[1][hirq] [12]),
        .I4(\slvo[3][hirq] [12]),
        .O(\slvi[hirq] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][12]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [12]),
        .I1(\msto[6][hirq] [12]),
        .I2(\msto[4][hirq] [12]),
        .I3(\msto[5][hirq] [12]),
        .I4(\msto[3][hirq] [12]),
        .I5(\msto[2][hirq] [12]),
        .O(\slvi[hirq][12]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][12]_INST_0_i_2 
       (.I0(\msto[0][hirq] [12]),
        .I1(\msto[1][hirq] [12]),
        .I2(\slvo[6][hirq] [12]),
        .I3(\slvo[7][hirq] [12]),
        .I4(\slvo[5][hirq] [12]),
        .I5(\slvo[4][hirq] [12]),
        .O(\slvi[hirq][12]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][13]_INST_0 
       (.I0(\slvi[hirq][13]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][13]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [13]),
        .I3(\slvo[1][hirq] [13]),
        .I4(\slvo[3][hirq] [13]),
        .O(\slvi[hirq] [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][13]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [13]),
        .I1(\msto[6][hirq] [13]),
        .I2(\msto[4][hirq] [13]),
        .I3(\msto[5][hirq] [13]),
        .I4(\msto[3][hirq] [13]),
        .I5(\msto[2][hirq] [13]),
        .O(\slvi[hirq][13]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][13]_INST_0_i_2 
       (.I0(\msto[0][hirq] [13]),
        .I1(\msto[1][hirq] [13]),
        .I2(\slvo[6][hirq] [13]),
        .I3(\slvo[7][hirq] [13]),
        .I4(\slvo[5][hirq] [13]),
        .I5(\slvo[4][hirq] [13]),
        .O(\slvi[hirq][13]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][14]_INST_0 
       (.I0(\slvi[hirq][14]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][14]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [14]),
        .I3(\slvo[1][hirq] [14]),
        .I4(\slvo[3][hirq] [14]),
        .O(\slvi[hirq] [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][14]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [14]),
        .I1(\msto[6][hirq] [14]),
        .I2(\msto[4][hirq] [14]),
        .I3(\msto[5][hirq] [14]),
        .I4(\msto[3][hirq] [14]),
        .I5(\msto[2][hirq] [14]),
        .O(\slvi[hirq][14]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][14]_INST_0_i_2 
       (.I0(\msto[0][hirq] [14]),
        .I1(\msto[1][hirq] [14]),
        .I2(\slvo[6][hirq] [14]),
        .I3(\slvo[7][hirq] [14]),
        .I4(\slvo[5][hirq] [14]),
        .I5(\slvo[4][hirq] [14]),
        .O(\slvi[hirq][14]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][15]_INST_0 
       (.I0(\slvi[hirq][15]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][15]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [15]),
        .I3(\slvo[1][hirq] [15]),
        .I4(\slvo[3][hirq] [15]),
        .O(\slvi[hirq] [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][15]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [15]),
        .I1(\msto[6][hirq] [15]),
        .I2(\msto[4][hirq] [15]),
        .I3(\msto[5][hirq] [15]),
        .I4(\msto[3][hirq] [15]),
        .I5(\msto[2][hirq] [15]),
        .O(\slvi[hirq][15]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][15]_INST_0_i_2 
       (.I0(\msto[0][hirq] [15]),
        .I1(\msto[1][hirq] [15]),
        .I2(\slvo[6][hirq] [15]),
        .I3(\slvo[7][hirq] [15]),
        .I4(\slvo[5][hirq] [15]),
        .I5(\slvo[4][hirq] [15]),
        .O(\slvi[hirq][15]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][16]_INST_0 
       (.I0(\slvi[hirq][16]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][16]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [16]),
        .I3(\slvo[1][hirq] [16]),
        .I4(\slvo[3][hirq] [16]),
        .O(\slvi[hirq] [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][16]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [16]),
        .I1(\msto[6][hirq] [16]),
        .I2(\msto[4][hirq] [16]),
        .I3(\msto[5][hirq] [16]),
        .I4(\msto[3][hirq] [16]),
        .I5(\msto[2][hirq] [16]),
        .O(\slvi[hirq][16]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][16]_INST_0_i_2 
       (.I0(\msto[0][hirq] [16]),
        .I1(\msto[1][hirq] [16]),
        .I2(\slvo[6][hirq] [16]),
        .I3(\slvo[7][hirq] [16]),
        .I4(\slvo[5][hirq] [16]),
        .I5(\slvo[4][hirq] [16]),
        .O(\slvi[hirq][16]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][17]_INST_0 
       (.I0(\slvi[hirq][17]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][17]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [17]),
        .I3(\slvo[1][hirq] [17]),
        .I4(\slvo[3][hirq] [17]),
        .O(\slvi[hirq] [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][17]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [17]),
        .I1(\msto[6][hirq] [17]),
        .I2(\msto[4][hirq] [17]),
        .I3(\msto[5][hirq] [17]),
        .I4(\msto[3][hirq] [17]),
        .I5(\msto[2][hirq] [17]),
        .O(\slvi[hirq][17]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][17]_INST_0_i_2 
       (.I0(\msto[0][hirq] [17]),
        .I1(\msto[1][hirq] [17]),
        .I2(\slvo[6][hirq] [17]),
        .I3(\slvo[7][hirq] [17]),
        .I4(\slvo[5][hirq] [17]),
        .I5(\slvo[4][hirq] [17]),
        .O(\slvi[hirq][17]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][18]_INST_0 
       (.I0(\slvi[hirq][18]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][18]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [18]),
        .I3(\slvo[1][hirq] [18]),
        .I4(\slvo[3][hirq] [18]),
        .O(\slvi[hirq] [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][18]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [18]),
        .I1(\msto[6][hirq] [18]),
        .I2(\msto[4][hirq] [18]),
        .I3(\msto[5][hirq] [18]),
        .I4(\msto[3][hirq] [18]),
        .I5(\msto[2][hirq] [18]),
        .O(\slvi[hirq][18]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][18]_INST_0_i_2 
       (.I0(\msto[0][hirq] [18]),
        .I1(\msto[1][hirq] [18]),
        .I2(\slvo[6][hirq] [18]),
        .I3(\slvo[7][hirq] [18]),
        .I4(\slvo[5][hirq] [18]),
        .I5(\slvo[4][hirq] [18]),
        .O(\slvi[hirq][18]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][19]_INST_0 
       (.I0(\slvi[hirq][19]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][19]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [19]),
        .I3(\slvo[1][hirq] [19]),
        .I4(\slvo[3][hirq] [19]),
        .O(\slvi[hirq] [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][19]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [19]),
        .I1(\msto[6][hirq] [19]),
        .I2(\msto[4][hirq] [19]),
        .I3(\msto[5][hirq] [19]),
        .I4(\msto[3][hirq] [19]),
        .I5(\msto[2][hirq] [19]),
        .O(\slvi[hirq][19]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][19]_INST_0_i_2 
       (.I0(\msto[0][hirq] [19]),
        .I1(\msto[1][hirq] [19]),
        .I2(\slvo[6][hirq] [19]),
        .I3(\slvo[7][hirq] [19]),
        .I4(\slvo[5][hirq] [19]),
        .I5(\slvo[4][hirq] [19]),
        .O(\slvi[hirq][19]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][1]_INST_0 
       (.I0(\slvi[hirq][1]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][1]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [1]),
        .I3(\slvo[1][hirq] [1]),
        .I4(\slvo[3][hirq] [1]),
        .O(\slvi[hirq] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][1]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [1]),
        .I1(\msto[6][hirq] [1]),
        .I2(\msto[4][hirq] [1]),
        .I3(\msto[5][hirq] [1]),
        .I4(\msto[3][hirq] [1]),
        .I5(\msto[2][hirq] [1]),
        .O(\slvi[hirq][1]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][1]_INST_0_i_2 
       (.I0(\msto[0][hirq] [1]),
        .I1(\msto[1][hirq] [1]),
        .I2(\slvo[6][hirq] [1]),
        .I3(\slvo[7][hirq] [1]),
        .I4(\slvo[5][hirq] [1]),
        .I5(\slvo[4][hirq] [1]),
        .O(\slvi[hirq][1]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][20]_INST_0 
       (.I0(\slvi[hirq][20]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][20]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [20]),
        .I3(\slvo[1][hirq] [20]),
        .I4(\slvo[3][hirq] [20]),
        .O(\slvi[hirq] [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][20]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [20]),
        .I1(\msto[6][hirq] [20]),
        .I2(\msto[4][hirq] [20]),
        .I3(\msto[5][hirq] [20]),
        .I4(\msto[3][hirq] [20]),
        .I5(\msto[2][hirq] [20]),
        .O(\slvi[hirq][20]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][20]_INST_0_i_2 
       (.I0(\msto[0][hirq] [20]),
        .I1(\msto[1][hirq] [20]),
        .I2(\slvo[6][hirq] [20]),
        .I3(\slvo[7][hirq] [20]),
        .I4(\slvo[5][hirq] [20]),
        .I5(\slvo[4][hirq] [20]),
        .O(\slvi[hirq][20]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][21]_INST_0 
       (.I0(\slvi[hirq][21]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][21]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [21]),
        .I3(\slvo[1][hirq] [21]),
        .I4(\slvo[3][hirq] [21]),
        .O(\slvi[hirq] [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][21]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [21]),
        .I1(\msto[6][hirq] [21]),
        .I2(\msto[4][hirq] [21]),
        .I3(\msto[5][hirq] [21]),
        .I4(\msto[3][hirq] [21]),
        .I5(\msto[2][hirq] [21]),
        .O(\slvi[hirq][21]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][21]_INST_0_i_2 
       (.I0(\msto[0][hirq] [21]),
        .I1(\msto[1][hirq] [21]),
        .I2(\slvo[6][hirq] [21]),
        .I3(\slvo[7][hirq] [21]),
        .I4(\slvo[5][hirq] [21]),
        .I5(\slvo[4][hirq] [21]),
        .O(\slvi[hirq][21]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][22]_INST_0 
       (.I0(\slvi[hirq][22]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][22]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [22]),
        .I3(\slvo[1][hirq] [22]),
        .I4(\slvo[3][hirq] [22]),
        .O(\slvi[hirq] [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][22]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [22]),
        .I1(\msto[6][hirq] [22]),
        .I2(\msto[4][hirq] [22]),
        .I3(\msto[5][hirq] [22]),
        .I4(\msto[3][hirq] [22]),
        .I5(\msto[2][hirq] [22]),
        .O(\slvi[hirq][22]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][22]_INST_0_i_2 
       (.I0(\msto[0][hirq] [22]),
        .I1(\msto[1][hirq] [22]),
        .I2(\slvo[6][hirq] [22]),
        .I3(\slvo[7][hirq] [22]),
        .I4(\slvo[5][hirq] [22]),
        .I5(\slvo[4][hirq] [22]),
        .O(\slvi[hirq][22]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][23]_INST_0 
       (.I0(\slvi[hirq][23]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][23]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [23]),
        .I3(\slvo[1][hirq] [23]),
        .I4(\slvo[3][hirq] [23]),
        .O(\slvi[hirq] [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][23]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [23]),
        .I1(\msto[6][hirq] [23]),
        .I2(\msto[4][hirq] [23]),
        .I3(\msto[5][hirq] [23]),
        .I4(\msto[3][hirq] [23]),
        .I5(\msto[2][hirq] [23]),
        .O(\slvi[hirq][23]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][23]_INST_0_i_2 
       (.I0(\msto[0][hirq] [23]),
        .I1(\msto[1][hirq] [23]),
        .I2(\slvo[6][hirq] [23]),
        .I3(\slvo[7][hirq] [23]),
        .I4(\slvo[5][hirq] [23]),
        .I5(\slvo[4][hirq] [23]),
        .O(\slvi[hirq][23]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][24]_INST_0 
       (.I0(\slvi[hirq][24]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][24]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [24]),
        .I3(\slvo[1][hirq] [24]),
        .I4(\slvo[3][hirq] [24]),
        .O(\slvi[hirq] [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][24]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [24]),
        .I1(\msto[6][hirq] [24]),
        .I2(\msto[4][hirq] [24]),
        .I3(\msto[5][hirq] [24]),
        .I4(\msto[3][hirq] [24]),
        .I5(\msto[2][hirq] [24]),
        .O(\slvi[hirq][24]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][24]_INST_0_i_2 
       (.I0(\msto[0][hirq] [24]),
        .I1(\msto[1][hirq] [24]),
        .I2(\slvo[6][hirq] [24]),
        .I3(\slvo[7][hirq] [24]),
        .I4(\slvo[5][hirq] [24]),
        .I5(\slvo[4][hirq] [24]),
        .O(\slvi[hirq][24]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][25]_INST_0 
       (.I0(\slvi[hirq][25]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][25]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [25]),
        .I3(\slvo[1][hirq] [25]),
        .I4(\slvo[3][hirq] [25]),
        .O(\slvi[hirq] [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][25]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [25]),
        .I1(\msto[6][hirq] [25]),
        .I2(\msto[4][hirq] [25]),
        .I3(\msto[5][hirq] [25]),
        .I4(\msto[3][hirq] [25]),
        .I5(\msto[2][hirq] [25]),
        .O(\slvi[hirq][25]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][25]_INST_0_i_2 
       (.I0(\msto[0][hirq] [25]),
        .I1(\msto[1][hirq] [25]),
        .I2(\slvo[6][hirq] [25]),
        .I3(\slvo[7][hirq] [25]),
        .I4(\slvo[5][hirq] [25]),
        .I5(\slvo[4][hirq] [25]),
        .O(\slvi[hirq][25]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][26]_INST_0 
       (.I0(\slvi[hirq][26]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][26]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [26]),
        .I3(\slvo[1][hirq] [26]),
        .I4(\slvo[3][hirq] [26]),
        .O(\slvi[hirq] [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][26]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [26]),
        .I1(\msto[6][hirq] [26]),
        .I2(\msto[4][hirq] [26]),
        .I3(\msto[5][hirq] [26]),
        .I4(\msto[3][hirq] [26]),
        .I5(\msto[2][hirq] [26]),
        .O(\slvi[hirq][26]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][26]_INST_0_i_2 
       (.I0(\msto[0][hirq] [26]),
        .I1(\msto[1][hirq] [26]),
        .I2(\slvo[6][hirq] [26]),
        .I3(\slvo[7][hirq] [26]),
        .I4(\slvo[5][hirq] [26]),
        .I5(\slvo[4][hirq] [26]),
        .O(\slvi[hirq][26]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][27]_INST_0 
       (.I0(\slvi[hirq][27]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][27]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [27]),
        .I3(\slvo[1][hirq] [27]),
        .I4(\slvo[3][hirq] [27]),
        .O(\slvi[hirq] [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][27]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [27]),
        .I1(\msto[6][hirq] [27]),
        .I2(\msto[4][hirq] [27]),
        .I3(\msto[5][hirq] [27]),
        .I4(\msto[3][hirq] [27]),
        .I5(\msto[2][hirq] [27]),
        .O(\slvi[hirq][27]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][27]_INST_0_i_2 
       (.I0(\msto[0][hirq] [27]),
        .I1(\msto[1][hirq] [27]),
        .I2(\slvo[6][hirq] [27]),
        .I3(\slvo[7][hirq] [27]),
        .I4(\slvo[5][hirq] [27]),
        .I5(\slvo[4][hirq] [27]),
        .O(\slvi[hirq][27]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][28]_INST_0 
       (.I0(\slvi[hirq][28]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][28]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [28]),
        .I3(\slvo[1][hirq] [28]),
        .I4(\slvo[3][hirq] [28]),
        .O(\slvi[hirq] [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][28]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [28]),
        .I1(\msto[6][hirq] [28]),
        .I2(\msto[4][hirq] [28]),
        .I3(\msto[5][hirq] [28]),
        .I4(\msto[3][hirq] [28]),
        .I5(\msto[2][hirq] [28]),
        .O(\slvi[hirq][28]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][28]_INST_0_i_2 
       (.I0(\msto[0][hirq] [28]),
        .I1(\msto[1][hirq] [28]),
        .I2(\slvo[6][hirq] [28]),
        .I3(\slvo[7][hirq] [28]),
        .I4(\slvo[5][hirq] [28]),
        .I5(\slvo[4][hirq] [28]),
        .O(\slvi[hirq][28]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][29]_INST_0 
       (.I0(\slvi[hirq][29]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][29]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [29]),
        .I3(\slvo[1][hirq] [29]),
        .I4(\slvo[3][hirq] [29]),
        .O(\slvi[hirq] [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][29]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [29]),
        .I1(\msto[6][hirq] [29]),
        .I2(\msto[4][hirq] [29]),
        .I3(\msto[5][hirq] [29]),
        .I4(\msto[3][hirq] [29]),
        .I5(\msto[2][hirq] [29]),
        .O(\slvi[hirq][29]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][29]_INST_0_i_2 
       (.I0(\msto[0][hirq] [29]),
        .I1(\msto[1][hirq] [29]),
        .I2(\slvo[6][hirq] [29]),
        .I3(\slvo[7][hirq] [29]),
        .I4(\slvo[5][hirq] [29]),
        .I5(\slvo[4][hirq] [29]),
        .O(\slvi[hirq][29]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][2]_INST_0 
       (.I0(\slvi[hirq][2]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][2]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [2]),
        .I3(\slvo[1][hirq] [2]),
        .I4(\slvo[3][hirq] [2]),
        .O(\slvi[hirq] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][2]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [2]),
        .I1(\msto[6][hirq] [2]),
        .I2(\msto[4][hirq] [2]),
        .I3(\msto[5][hirq] [2]),
        .I4(\msto[3][hirq] [2]),
        .I5(\msto[2][hirq] [2]),
        .O(\slvi[hirq][2]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][2]_INST_0_i_2 
       (.I0(\msto[0][hirq] [2]),
        .I1(\msto[1][hirq] [2]),
        .I2(\slvo[6][hirq] [2]),
        .I3(\slvo[7][hirq] [2]),
        .I4(\slvo[5][hirq] [2]),
        .I5(\slvo[4][hirq] [2]),
        .O(\slvi[hirq][2]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][30]_INST_0 
       (.I0(\slvi[hirq][30]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][30]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [30]),
        .I3(\slvo[1][hirq] [30]),
        .I4(\slvo[3][hirq] [30]),
        .O(\slvi[hirq] [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][30]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [30]),
        .I1(\msto[6][hirq] [30]),
        .I2(\msto[4][hirq] [30]),
        .I3(\msto[5][hirq] [30]),
        .I4(\msto[3][hirq] [30]),
        .I5(\msto[2][hirq] [30]),
        .O(\slvi[hirq][30]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][30]_INST_0_i_2 
       (.I0(\msto[0][hirq] [30]),
        .I1(\msto[1][hirq] [30]),
        .I2(\slvo[6][hirq] [30]),
        .I3(\slvo[7][hirq] [30]),
        .I4(\slvo[5][hirq] [30]),
        .I5(\slvo[4][hirq] [30]),
        .O(\slvi[hirq][30]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][31]_INST_0 
       (.I0(\slvi[hirq][31]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][31]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [31]),
        .I3(\slvo[1][hirq] [31]),
        .I4(\slvo[3][hirq] [31]),
        .O(\slvi[hirq] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][31]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [31]),
        .I1(\msto[6][hirq] [31]),
        .I2(\msto[4][hirq] [31]),
        .I3(\msto[5][hirq] [31]),
        .I4(\msto[3][hirq] [31]),
        .I5(\msto[2][hirq] [31]),
        .O(\slvi[hirq][31]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][31]_INST_0_i_2 
       (.I0(\msto[0][hirq] [31]),
        .I1(\msto[1][hirq] [31]),
        .I2(\slvo[6][hirq] [31]),
        .I3(\slvo[7][hirq] [31]),
        .I4(\slvo[5][hirq] [31]),
        .I5(\slvo[4][hirq] [31]),
        .O(\slvi[hirq][31]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][3]_INST_0 
       (.I0(\slvi[hirq][3]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][3]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [3]),
        .I3(\slvo[1][hirq] [3]),
        .I4(\slvo[3][hirq] [3]),
        .O(\slvi[hirq] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][3]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [3]),
        .I1(\msto[6][hirq] [3]),
        .I2(\msto[4][hirq] [3]),
        .I3(\msto[5][hirq] [3]),
        .I4(\msto[3][hirq] [3]),
        .I5(\msto[2][hirq] [3]),
        .O(\slvi[hirq][3]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][3]_INST_0_i_2 
       (.I0(\msto[0][hirq] [3]),
        .I1(\msto[1][hirq] [3]),
        .I2(\slvo[6][hirq] [3]),
        .I3(\slvo[7][hirq] [3]),
        .I4(\slvo[5][hirq] [3]),
        .I5(\slvo[4][hirq] [3]),
        .O(\slvi[hirq][3]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][4]_INST_0 
       (.I0(\slvi[hirq][4]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][4]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [4]),
        .I3(\slvo[1][hirq] [4]),
        .I4(\slvo[3][hirq] [4]),
        .O(\slvi[hirq] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][4]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [4]),
        .I1(\msto[6][hirq] [4]),
        .I2(\msto[4][hirq] [4]),
        .I3(\msto[5][hirq] [4]),
        .I4(\msto[3][hirq] [4]),
        .I5(\msto[2][hirq] [4]),
        .O(\slvi[hirq][4]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][4]_INST_0_i_2 
       (.I0(\msto[0][hirq] [4]),
        .I1(\msto[1][hirq] [4]),
        .I2(\slvo[6][hirq] [4]),
        .I3(\slvo[7][hirq] [4]),
        .I4(\slvo[5][hirq] [4]),
        .I5(\slvo[4][hirq] [4]),
        .O(\slvi[hirq][4]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][5]_INST_0 
       (.I0(\slvi[hirq][5]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][5]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [5]),
        .I3(\slvo[1][hirq] [5]),
        .I4(\slvo[3][hirq] [5]),
        .O(\slvi[hirq] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][5]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [5]),
        .I1(\msto[6][hirq] [5]),
        .I2(\msto[4][hirq] [5]),
        .I3(\msto[5][hirq] [5]),
        .I4(\msto[3][hirq] [5]),
        .I5(\msto[2][hirq] [5]),
        .O(\slvi[hirq][5]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][5]_INST_0_i_2 
       (.I0(\msto[0][hirq] [5]),
        .I1(\msto[1][hirq] [5]),
        .I2(\slvo[6][hirq] [5]),
        .I3(\slvo[7][hirq] [5]),
        .I4(\slvo[5][hirq] [5]),
        .I5(\slvo[4][hirq] [5]),
        .O(\slvi[hirq][5]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][6]_INST_0 
       (.I0(\slvi[hirq][6]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][6]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [6]),
        .I3(\slvo[1][hirq] [6]),
        .I4(\slvo[3][hirq] [6]),
        .O(\slvi[hirq] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][6]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [6]),
        .I1(\msto[6][hirq] [6]),
        .I2(\msto[4][hirq] [6]),
        .I3(\msto[5][hirq] [6]),
        .I4(\msto[3][hirq] [6]),
        .I5(\msto[2][hirq] [6]),
        .O(\slvi[hirq][6]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][6]_INST_0_i_2 
       (.I0(\msto[0][hirq] [6]),
        .I1(\msto[1][hirq] [6]),
        .I2(\slvo[6][hirq] [6]),
        .I3(\slvo[7][hirq] [6]),
        .I4(\slvo[5][hirq] [6]),
        .I5(\slvo[4][hirq] [6]),
        .O(\slvi[hirq][6]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][7]_INST_0 
       (.I0(\slvi[hirq][7]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][7]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [7]),
        .I3(\slvo[1][hirq] [7]),
        .I4(\slvo[3][hirq] [7]),
        .O(\slvi[hirq] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][7]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [7]),
        .I1(\msto[6][hirq] [7]),
        .I2(\msto[4][hirq] [7]),
        .I3(\msto[5][hirq] [7]),
        .I4(\msto[3][hirq] [7]),
        .I5(\msto[2][hirq] [7]),
        .O(\slvi[hirq][7]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][7]_INST_0_i_2 
       (.I0(\msto[0][hirq] [7]),
        .I1(\msto[1][hirq] [7]),
        .I2(\slvo[6][hirq] [7]),
        .I3(\slvo[7][hirq] [7]),
        .I4(\slvo[5][hirq] [7]),
        .I5(\slvo[4][hirq] [7]),
        .O(\slvi[hirq][7]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][8]_INST_0 
       (.I0(\slvi[hirq][8]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][8]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [8]),
        .I3(\slvo[1][hirq] [8]),
        .I4(\slvo[3][hirq] [8]),
        .O(\slvi[hirq] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][8]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [8]),
        .I1(\msto[6][hirq] [8]),
        .I2(\msto[4][hirq] [8]),
        .I3(\msto[5][hirq] [8]),
        .I4(\msto[3][hirq] [8]),
        .I5(\msto[2][hirq] [8]),
        .O(\slvi[hirq][8]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][8]_INST_0_i_2 
       (.I0(\msto[0][hirq] [8]),
        .I1(\msto[1][hirq] [8]),
        .I2(\slvo[6][hirq] [8]),
        .I3(\slvo[7][hirq] [8]),
        .I4(\slvo[5][hirq] [8]),
        .I5(\slvo[4][hirq] [8]),
        .O(\slvi[hirq][8]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \slvi[hirq][9]_INST_0 
       (.I0(\slvi[hirq][9]_INST_0_i_1_n_0 ),
        .I1(\slvi[hirq][9]_INST_0_i_2_n_0 ),
        .I2(\slvo[2][hirq] [9]),
        .I3(\slvo[1][hirq] [9]),
        .I4(\slvo[3][hirq] [9]),
        .O(\slvi[hirq] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][9]_INST_0_i_1 
       (.I0(\slvo[0][hirq] [9]),
        .I1(\msto[6][hirq] [9]),
        .I2(\msto[4][hirq] [9]),
        .I3(\msto[5][hirq] [9]),
        .I4(\msto[3][hirq] [9]),
        .I5(\msto[2][hirq] [9]),
        .O(\slvi[hirq][9]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \slvi[hirq][9]_INST_0_i_2 
       (.I0(\msto[0][hirq] [9]),
        .I1(\msto[1][hirq] [9]),
        .I2(\slvo[6][hirq] [9]),
        .I3(\slvo[7][hirq] [9]),
        .I4(\slvo[5][hirq] [9]),
        .I5(\slvo[4][hirq] [9]),
        .O(\slvi[hirq][9]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF7FFFFFFFFFFFFFF)) 
    \slvi[hmbsel][0]_INST_0 
       (.I0(\slvi[hmbsel][0]_INST_0_i_1_n_0 ),
        .I1(\slvi[hmbsel][0]_INST_0_i_2_n_0 ),
        .I2(\slvi[hmbsel][0]_INST_0_i_3_n_0 ),
        .I3(\slvi[hmbsel][0]_INST_0_i_4_n_0 ),
        .I4(\slvi[hmbsel][0]_INST_0_i_5_n_0 ),
        .I5(\slvi[hmbsel][0]_INST_0_i_6_n_0 ),
        .O(\slvi[hmbsel] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][0]_INST_0_i_1 
       (.I0(\slvo[6][hconfig][4] [1]),
        .I1(\slvi[hmbsel][0]_INST_0_i_7_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \slvi[hmbsel][0]_INST_0_i_10 
       (.I0(hsel2168_in),
        .I1(hsel358_out),
        .I2(hsel219_in),
        .O(hsel1169_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_100 
       (.I0(\slvo[3][hconfig][4] [11]),
        .I1(\slvo[3][hconfig][4] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[3][hconfig][4] [12]),
        .I4(\slvo[3][hconfig][4] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hmbsel][0]_INST_0_i_100_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_101 
       (.I0(\slvo[3][hconfig][4] [8]),
        .I1(\slvo[3][hconfig][4] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[3][hconfig][4] [9]),
        .I4(\slvo[3][hconfig][4] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hmbsel][0]_INST_0_i_101_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_102 
       (.I0(\slvo[3][hconfig][4] [5]),
        .I1(\slvo[3][hconfig][4] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[3][hconfig][4] [6]),
        .I4(\slvo[3][hconfig][4] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hmbsel][0]_INST_0_i_102_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_103 
       (.I0(\slvo[5][hconfig][4] [14]),
        .I1(\slvo[5][hconfig][4] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[5][hconfig][4] [15]),
        .I4(\slvo[5][hconfig][4] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hmbsel][0]_INST_0_i_103_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_104 
       (.I0(\slvo[5][hconfig][4] [11]),
        .I1(\slvo[5][hconfig][4] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[5][hconfig][4] [12]),
        .I4(\slvo[5][hconfig][4] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hmbsel][0]_INST_0_i_104_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_105 
       (.I0(\slvo[5][hconfig][4] [8]),
        .I1(\slvo[5][hconfig][4] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[5][hconfig][4] [9]),
        .I4(\slvo[5][hconfig][4] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hmbsel][0]_INST_0_i_105_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_106 
       (.I0(\slvo[5][hconfig][4] [5]),
        .I1(\slvo[5][hconfig][4] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[5][hconfig][4] [6]),
        .I4(\slvo[5][hconfig][4] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hmbsel][0]_INST_0_i_106_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_107 
       (.I0(\slvo[5][hconfig][4] [14]),
        .I1(\slvo[5][hconfig][4] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[5][hconfig][4] [15]),
        .I4(\slvo[5][hconfig][4] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hmbsel][0]_INST_0_i_107_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_108 
       (.I0(\slvo[5][hconfig][4] [11]),
        .I1(\slvo[5][hconfig][4] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[5][hconfig][4] [12]),
        .I4(\slvo[5][hconfig][4] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hmbsel][0]_INST_0_i_108_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_109 
       (.I0(\slvo[5][hconfig][4] [8]),
        .I1(\slvo[5][hconfig][4] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[5][hconfig][4] [9]),
        .I4(\slvo[5][hconfig][4] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hmbsel][0]_INST_0_i_109_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000808030003000)) 
    \slvi[hmbsel][0]_INST_0_i_11 
       (.I0(hsel334_out),
        .I1(\slvo[3][hconfig][4] [0]),
        .I2(hsel2108_in),
        .I3(hsel335_out),
        .I4(\slvi[hmbsel][2]_INST_0_i_9_n_0 ),
        .I5(\slvi[hmbsel][2]_INST_0_i_10_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_110 
       (.I0(\slvo[5][hconfig][4] [5]),
        .I1(\slvo[5][hconfig][4] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[5][hconfig][4] [6]),
        .I4(\slvo[5][hconfig][4] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hmbsel][0]_INST_0_i_110_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_111 
       (.I0(\slvo[7][hconfig][4] [14]),
        .I1(\slvo[7][hconfig][4] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[7][hconfig][4] [15]),
        .I4(\slvo[7][hconfig][4] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hmbsel][0]_INST_0_i_111_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_112 
       (.I0(\slvo[7][hconfig][4] [11]),
        .I1(\slvo[7][hconfig][4] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[7][hconfig][4] [12]),
        .I4(\slvo[7][hconfig][4] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hmbsel][0]_INST_0_i_112_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_113 
       (.I0(\slvo[7][hconfig][4] [8]),
        .I1(\slvo[7][hconfig][4] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[7][hconfig][4] [9]),
        .I4(\slvo[7][hconfig][4] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hmbsel][0]_INST_0_i_113_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_114 
       (.I0(\slvo[7][hconfig][4] [5]),
        .I1(\slvo[7][hconfig][4] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[7][hconfig][4] [6]),
        .I4(\slvo[7][hconfig][4] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hmbsel][0]_INST_0_i_114_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_115 
       (.I0(\slvo[7][hconfig][4] [14]),
        .I1(\slvo[7][hconfig][4] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[7][hconfig][4] [15]),
        .I4(\slvo[7][hconfig][4] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hmbsel][0]_INST_0_i_115_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_116 
       (.I0(\slvo[7][hconfig][4] [11]),
        .I1(\slvo[7][hconfig][4] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[7][hconfig][4] [12]),
        .I4(\slvo[7][hconfig][4] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hmbsel][0]_INST_0_i_116_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_117 
       (.I0(\slvo[7][hconfig][4] [8]),
        .I1(\slvo[7][hconfig][4] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[7][hconfig][4] [9]),
        .I4(\slvo[7][hconfig][4] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hmbsel][0]_INST_0_i_117_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_118 
       (.I0(\slvo[7][hconfig][4] [5]),
        .I1(\slvo[7][hconfig][4] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[7][hconfig][4] [6]),
        .I4(\slvo[7][hconfig][4] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hmbsel][0]_INST_0_i_118_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000808030003000)) 
    \slvi[hmbsel][0]_INST_0_i_12 
       (.I0(hsel318_out),
        .I1(\slvo[5][hconfig][4] [0]),
        .I2(hsel268_in),
        .I3(hsel319_out),
        .I4(\slvi[hmbsel][2]_INST_0_i_9_n_0 ),
        .I5(\slvi[hmbsel][2]_INST_0_i_10_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000808030003000)) 
    \slvi[hmbsel][0]_INST_0_i_13 
       (.I0(hsel32_out),
        .I1(\slvo[7][hconfig][4] [0]),
        .I2(hsel227_in),
        .I3(hsel33_out),
        .I4(\slvi[hmbsel][2]_INST_0_i_9_n_0 ),
        .I5(\slvi[hmbsel][2]_INST_0_i_10_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][0]_INST_0_i_14 
       (.CI(slvi),
        .CO({hsel310_out,\slvi[hmbsel][0]_INST_0_i_14_n_1 ,\slvi[hmbsel][0]_INST_0_i_14_n_2 ,\slvi[hmbsel][0]_INST_0_i_14_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][0]_INST_0_i_29_n_0 ,\slvi[hmbsel][0]_INST_0_i_30_n_0 ,\slvi[hmbsel][0]_INST_0_i_31_n_0 ,\slvi[hmbsel][0]_INST_0_i_32_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][0]_INST_0_i_15 
       (.I0(\slvi[hmbsel][0]_INST_0_i_33_n_0 ),
        .I1(\slvi[hmbsel][0]_INST_0_i_34_n_0 ),
        .O(hsel248_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][0]_INST_0_i_16 
       (.CI(slvi),
        .CO({hsel311_out,\slvi[hmbsel][0]_INST_0_i_16_n_1 ,\slvi[hmbsel][0]_INST_0_i_16_n_2 ,\slvi[hmbsel][0]_INST_0_i_16_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][0]_INST_0_i_35_n_0 ,\slvi[hmbsel][0]_INST_0_i_36_n_0 ,\slvi[hmbsel][0]_INST_0_i_37_n_0 ,\slvi[hmbsel][0]_INST_0_i_38_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][0]_INST_0_i_17 
       (.CI(slvi),
        .CO({hsel326_out,\slvi[hmbsel][0]_INST_0_i_17_n_1 ,\slvi[hmbsel][0]_INST_0_i_17_n_2 ,\slvi[hmbsel][0]_INST_0_i_17_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][0]_INST_0_i_39_n_0 ,\slvi[hmbsel][0]_INST_0_i_40_n_0 ,\slvi[hmbsel][0]_INST_0_i_41_n_0 ,\slvi[hmbsel][0]_INST_0_i_42_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][0]_INST_0_i_18 
       (.I0(\slvi[hmbsel][0]_INST_0_i_43_n_0 ),
        .I1(\slvi[hmbsel][0]_INST_0_i_44_n_0 ),
        .O(hsel288_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][0]_INST_0_i_19 
       (.CI(slvi),
        .CO({hsel327_out,\slvi[hmbsel][0]_INST_0_i_19_n_1 ,\slvi[hmbsel][0]_INST_0_i_19_n_2 ,\slvi[hmbsel][0]_INST_0_i_19_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][0]_INST_0_i_45_n_0 ,\slvi[hmbsel][0]_INST_0_i_46_n_0 ,\slvi[hmbsel][0]_INST_0_i_47_n_0 ,\slvi[hmbsel][0]_INST_0_i_48_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][0]_INST_0_i_2 
       (.I0(\slvo[4][hconfig][4] [1]),
        .I1(\slvi[hmbsel][0]_INST_0_i_8_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][0]_INST_0_i_20 
       (.CI(slvi),
        .CO({hsel334_out,\slvi[hmbsel][0]_INST_0_i_20_n_1 ,\slvi[hmbsel][0]_INST_0_i_20_n_2 ,\slvi[hmbsel][0]_INST_0_i_20_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][0]_INST_0_i_49_n_0 ,\slvi[hmbsel][0]_INST_0_i_50_n_0 ,\slvi[hmbsel][0]_INST_0_i_51_n_0 ,\slvi[hmbsel][0]_INST_0_i_52_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][0]_INST_0_i_21 
       (.I0(\slvi[hmbsel][0]_INST_0_i_53_n_0 ),
        .I1(\slvi[hmbsel][0]_INST_0_i_54_n_0 ),
        .O(hsel2108_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][0]_INST_0_i_22 
       (.CI(slvi),
        .CO({hsel335_out,\slvi[hmbsel][0]_INST_0_i_22_n_1 ,\slvi[hmbsel][0]_INST_0_i_22_n_2 ,\slvi[hmbsel][0]_INST_0_i_22_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][0]_INST_0_i_55_n_0 ,\slvi[hmbsel][0]_INST_0_i_56_n_0 ,\slvi[hmbsel][0]_INST_0_i_57_n_0 ,\slvi[hmbsel][0]_INST_0_i_58_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][0]_INST_0_i_23 
       (.CI(slvi),
        .CO({hsel318_out,\slvi[hmbsel][0]_INST_0_i_23_n_1 ,\slvi[hmbsel][0]_INST_0_i_23_n_2 ,\slvi[hmbsel][0]_INST_0_i_23_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][0]_INST_0_i_59_n_0 ,\slvi[hmbsel][0]_INST_0_i_60_n_0 ,\slvi[hmbsel][0]_INST_0_i_61_n_0 ,\slvi[hmbsel][0]_INST_0_i_62_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][0]_INST_0_i_24 
       (.I0(\slvi[hmbsel][0]_INST_0_i_63_n_0 ),
        .I1(\slvi[hmbsel][0]_INST_0_i_64_n_0 ),
        .O(hsel268_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][0]_INST_0_i_25 
       (.CI(slvi),
        .CO({hsel319_out,\slvi[hmbsel][0]_INST_0_i_25_n_1 ,\slvi[hmbsel][0]_INST_0_i_25_n_2 ,\slvi[hmbsel][0]_INST_0_i_25_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][0]_INST_0_i_65_n_0 ,\slvi[hmbsel][0]_INST_0_i_66_n_0 ,\slvi[hmbsel][0]_INST_0_i_67_n_0 ,\slvi[hmbsel][0]_INST_0_i_68_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][0]_INST_0_i_26 
       (.CI(slvi),
        .CO({hsel32_out,\slvi[hmbsel][0]_INST_0_i_26_n_1 ,\slvi[hmbsel][0]_INST_0_i_26_n_2 ,\slvi[hmbsel][0]_INST_0_i_26_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][0]_INST_0_i_69_n_0 ,\slvi[hmbsel][0]_INST_0_i_70_n_0 ,\slvi[hmbsel][0]_INST_0_i_71_n_0 ,\slvi[hmbsel][0]_INST_0_i_72_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][0]_INST_0_i_27 
       (.I0(\slvi[hmbsel][0]_INST_0_i_73_n_0 ),
        .I1(\slvi[hmbsel][0]_INST_0_i_74_n_0 ),
        .O(hsel227_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][0]_INST_0_i_28 
       (.CI(slvi),
        .CO({hsel33_out,\slvi[hmbsel][0]_INST_0_i_28_n_1 ,\slvi[hmbsel][0]_INST_0_i_28_n_2 ,\slvi[hmbsel][0]_INST_0_i_28_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][0]_INST_0_i_75_n_0 ,\slvi[hmbsel][0]_INST_0_i_76_n_0 ,\slvi[hmbsel][0]_INST_0_i_77_n_0 ,\slvi[hmbsel][0]_INST_0_i_78_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_29 
       (.I0(\slvo[6][hconfig][4] [13]),
        .I1(\slvo[6][hconfig][4] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hmbsel][0]_INST_0_i_79_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDD555D5FFFFFFFF)) 
    \slvi[hmbsel][0]_INST_0_i_3 
       (.I0(\slvi[hsel][1]_INST_0_i_2_n_0 ),
        .I1(\slvo[0][hconfig][4] [1]),
        .I2(hsel1171_out),
        .I3(\slvo[0][hconfig][4] [0]),
        .I4(hsel1169_out),
        .I5(\slvi[hsel][2]_INST_0_i_3_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_30 
       (.I0(\slvo[6][hconfig][4] [10]),
        .I1(\slvo[6][hconfig][4] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hmbsel][0]_INST_0_i_80_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_31 
       (.I0(\slvo[6][hconfig][4] [7]),
        .I1(\slvo[6][hconfig][4] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hmbsel][0]_INST_0_i_81_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_32 
       (.I0(\slvo[6][hconfig][4] [4]),
        .I1(\slvo[6][hconfig][4] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hmbsel][0]_INST_0_i_82_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][0]_INST_0_i_33 
       (.I0(\slvo[6][hconfig][4] [9]),
        .I1(\slvo[6][hconfig][4] [7]),
        .I2(\slvo[6][hconfig][4] [8]),
        .I3(\slvo[6][hconfig][4] [4]),
        .I4(\slvo[6][hconfig][4] [5]),
        .I5(\slvo[6][hconfig][4] [6]),
        .O(\slvi[hmbsel][0]_INST_0_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][0]_INST_0_i_34 
       (.I0(\slvo[6][hconfig][4] [14]),
        .I1(\slvo[6][hconfig][4] [13]),
        .I2(\slvo[6][hconfig][4] [15]),
        .I3(\slvo[6][hconfig][4] [10]),
        .I4(\slvo[6][hconfig][4] [11]),
        .I5(\slvo[6][hconfig][4] [12]),
        .O(\slvi[hmbsel][0]_INST_0_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_35 
       (.I0(\slvo[6][hconfig][4] [13]),
        .I1(\slvo[6][hconfig][4] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hmbsel][0]_INST_0_i_83_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_36 
       (.I0(\slvo[6][hconfig][4] [10]),
        .I1(\slvo[6][hconfig][4] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hmbsel][0]_INST_0_i_84_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_37 
       (.I0(\slvo[6][hconfig][4] [7]),
        .I1(\slvo[6][hconfig][4] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hmbsel][0]_INST_0_i_85_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_38 
       (.I0(\slvo[6][hconfig][4] [4]),
        .I1(\slvo[6][hconfig][4] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hmbsel][0]_INST_0_i_86_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_39 
       (.I0(\slvo[4][hconfig][4] [13]),
        .I1(\slvo[4][hconfig][4] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hmbsel][0]_INST_0_i_87_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][0]_INST_0_i_4 
       (.I0(\slvo[3][hconfig][4] [1]),
        .I1(\slvi[hmbsel][0]_INST_0_i_11_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_40 
       (.I0(\slvo[4][hconfig][4] [10]),
        .I1(\slvo[4][hconfig][4] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hmbsel][0]_INST_0_i_88_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_41 
       (.I0(\slvo[4][hconfig][4] [7]),
        .I1(\slvo[4][hconfig][4] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hmbsel][0]_INST_0_i_89_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_42 
       (.I0(\slvo[4][hconfig][4] [4]),
        .I1(\slvo[4][hconfig][4] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hmbsel][0]_INST_0_i_90_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][0]_INST_0_i_43 
       (.I0(\slvo[4][hconfig][4] [9]),
        .I1(\slvo[4][hconfig][4] [7]),
        .I2(\slvo[4][hconfig][4] [8]),
        .I3(\slvo[4][hconfig][4] [4]),
        .I4(\slvo[4][hconfig][4] [5]),
        .I5(\slvo[4][hconfig][4] [6]),
        .O(\slvi[hmbsel][0]_INST_0_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][0]_INST_0_i_44 
       (.I0(\slvo[4][hconfig][4] [14]),
        .I1(\slvo[4][hconfig][4] [13]),
        .I2(\slvo[4][hconfig][4] [15]),
        .I3(\slvo[4][hconfig][4] [10]),
        .I4(\slvo[4][hconfig][4] [11]),
        .I5(\slvo[4][hconfig][4] [12]),
        .O(\slvi[hmbsel][0]_INST_0_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_45 
       (.I0(\slvo[4][hconfig][4] [13]),
        .I1(\slvo[4][hconfig][4] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hmbsel][0]_INST_0_i_91_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_46 
       (.I0(\slvo[4][hconfig][4] [10]),
        .I1(\slvo[4][hconfig][4] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hmbsel][0]_INST_0_i_92_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_47 
       (.I0(\slvo[4][hconfig][4] [7]),
        .I1(\slvo[4][hconfig][4] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hmbsel][0]_INST_0_i_93_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_48 
       (.I0(\slvo[4][hconfig][4] [4]),
        .I1(\slvo[4][hconfig][4] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hmbsel][0]_INST_0_i_94_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_49 
       (.I0(\slvo[3][hconfig][4] [13]),
        .I1(\slvo[3][hconfig][4] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hmbsel][0]_INST_0_i_95_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][0]_INST_0_i_5 
       (.I0(\slvo[5][hconfig][4] [1]),
        .I1(\slvi[hmbsel][0]_INST_0_i_12_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_50 
       (.I0(\slvo[3][hconfig][4] [10]),
        .I1(\slvo[3][hconfig][4] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hmbsel][0]_INST_0_i_96_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_51 
       (.I0(\slvo[3][hconfig][4] [7]),
        .I1(\slvo[3][hconfig][4] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hmbsel][0]_INST_0_i_97_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_51_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_52 
       (.I0(\slvo[3][hconfig][4] [4]),
        .I1(\slvo[3][hconfig][4] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hmbsel][0]_INST_0_i_98_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_52_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][0]_INST_0_i_53 
       (.I0(\slvo[3][hconfig][4] [9]),
        .I1(\slvo[3][hconfig][4] [7]),
        .I2(\slvo[3][hconfig][4] [8]),
        .I3(\slvo[3][hconfig][4] [4]),
        .I4(\slvo[3][hconfig][4] [5]),
        .I5(\slvo[3][hconfig][4] [6]),
        .O(\slvi[hmbsel][0]_INST_0_i_53_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][0]_INST_0_i_54 
       (.I0(\slvo[3][hconfig][4] [14]),
        .I1(\slvo[3][hconfig][4] [13]),
        .I2(\slvo[3][hconfig][4] [15]),
        .I3(\slvo[3][hconfig][4] [10]),
        .I4(\slvo[3][hconfig][4] [11]),
        .I5(\slvo[3][hconfig][4] [12]),
        .O(\slvi[hmbsel][0]_INST_0_i_54_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_55 
       (.I0(\slvo[3][hconfig][4] [13]),
        .I1(\slvo[3][hconfig][4] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hmbsel][0]_INST_0_i_99_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_55_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_56 
       (.I0(\slvo[3][hconfig][4] [10]),
        .I1(\slvo[3][hconfig][4] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hmbsel][0]_INST_0_i_100_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_56_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_57 
       (.I0(\slvo[3][hconfig][4] [7]),
        .I1(\slvo[3][hconfig][4] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hmbsel][0]_INST_0_i_101_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_57_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_58 
       (.I0(\slvo[3][hconfig][4] [4]),
        .I1(\slvo[3][hconfig][4] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hmbsel][0]_INST_0_i_102_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_58_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_59 
       (.I0(\slvo[5][hconfig][4] [13]),
        .I1(\slvo[5][hconfig][4] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hmbsel][0]_INST_0_i_103_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_59_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][0]_INST_0_i_6 
       (.I0(\slvo[7][hconfig][4] [1]),
        .I1(\slvi[hmbsel][0]_INST_0_i_13_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_60 
       (.I0(\slvo[5][hconfig][4] [10]),
        .I1(\slvo[5][hconfig][4] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hmbsel][0]_INST_0_i_104_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_60_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_61 
       (.I0(\slvo[5][hconfig][4] [7]),
        .I1(\slvo[5][hconfig][4] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hmbsel][0]_INST_0_i_105_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_61_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_62 
       (.I0(\slvo[5][hconfig][4] [4]),
        .I1(\slvo[5][hconfig][4] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hmbsel][0]_INST_0_i_106_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_62_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][0]_INST_0_i_63 
       (.I0(\slvo[5][hconfig][4] [9]),
        .I1(\slvo[5][hconfig][4] [7]),
        .I2(\slvo[5][hconfig][4] [8]),
        .I3(\slvo[5][hconfig][4] [4]),
        .I4(\slvo[5][hconfig][4] [5]),
        .I5(\slvo[5][hconfig][4] [6]),
        .O(\slvi[hmbsel][0]_INST_0_i_63_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][0]_INST_0_i_64 
       (.I0(\slvo[5][hconfig][4] [14]),
        .I1(\slvo[5][hconfig][4] [13]),
        .I2(\slvo[5][hconfig][4] [15]),
        .I3(\slvo[5][hconfig][4] [10]),
        .I4(\slvo[5][hconfig][4] [11]),
        .I5(\slvo[5][hconfig][4] [12]),
        .O(\slvi[hmbsel][0]_INST_0_i_64_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_65 
       (.I0(\slvo[5][hconfig][4] [13]),
        .I1(\slvo[5][hconfig][4] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hmbsel][0]_INST_0_i_107_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_65_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_66 
       (.I0(\slvo[5][hconfig][4] [10]),
        .I1(\slvo[5][hconfig][4] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hmbsel][0]_INST_0_i_108_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_66_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_67 
       (.I0(\slvo[5][hconfig][4] [7]),
        .I1(\slvo[5][hconfig][4] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hmbsel][0]_INST_0_i_109_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_67_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_68 
       (.I0(\slvo[5][hconfig][4] [4]),
        .I1(\slvo[5][hconfig][4] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hmbsel][0]_INST_0_i_110_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_68_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_69 
       (.I0(\slvo[7][hconfig][4] [13]),
        .I1(\slvo[7][hconfig][4] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hmbsel][0]_INST_0_i_111_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_69_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000808030003000)) 
    \slvi[hmbsel][0]_INST_0_i_7 
       (.I0(hsel310_out),
        .I1(\slvo[6][hconfig][4] [0]),
        .I2(hsel248_in),
        .I3(hsel311_out),
        .I4(\slvi[hmbsel][2]_INST_0_i_9_n_0 ),
        .I5(\slvi[hmbsel][2]_INST_0_i_10_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_70 
       (.I0(\slvo[7][hconfig][4] [10]),
        .I1(\slvo[7][hconfig][4] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hmbsel][0]_INST_0_i_112_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_70_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_71 
       (.I0(\slvo[7][hconfig][4] [7]),
        .I1(\slvo[7][hconfig][4] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hmbsel][0]_INST_0_i_113_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_71_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_72 
       (.I0(\slvo[7][hconfig][4] [4]),
        .I1(\slvo[7][hconfig][4] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hmbsel][0]_INST_0_i_114_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_72_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][0]_INST_0_i_73 
       (.I0(\slvo[7][hconfig][4] [9]),
        .I1(\slvo[7][hconfig][4] [7]),
        .I2(\slvo[7][hconfig][4] [8]),
        .I3(\slvo[7][hconfig][4] [4]),
        .I4(\slvo[7][hconfig][4] [5]),
        .I5(\slvo[7][hconfig][4] [6]),
        .O(\slvi[hmbsel][0]_INST_0_i_73_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][0]_INST_0_i_74 
       (.I0(\slvo[7][hconfig][4] [14]),
        .I1(\slvo[7][hconfig][4] [13]),
        .I2(\slvo[7][hconfig][4] [15]),
        .I3(\slvo[7][hconfig][4] [10]),
        .I4(\slvo[7][hconfig][4] [11]),
        .I5(\slvo[7][hconfig][4] [12]),
        .O(\slvi[hmbsel][0]_INST_0_i_74_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_75 
       (.I0(\slvo[7][hconfig][4] [13]),
        .I1(\slvo[7][hconfig][4] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hmbsel][0]_INST_0_i_115_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_75_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_76 
       (.I0(\slvo[7][hconfig][4] [10]),
        .I1(\slvo[7][hconfig][4] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hmbsel][0]_INST_0_i_116_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_76_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_77 
       (.I0(\slvo[7][hconfig][4] [7]),
        .I1(\slvo[7][hconfig][4] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hmbsel][0]_INST_0_i_117_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_77_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][0]_INST_0_i_78 
       (.I0(\slvo[7][hconfig][4] [4]),
        .I1(\slvo[7][hconfig][4] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hmbsel][0]_INST_0_i_118_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_78_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_79 
       (.I0(\slvo[6][hconfig][4] [14]),
        .I1(\slvo[6][hconfig][4] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[6][hconfig][4] [15]),
        .I4(\slvo[6][hconfig][4] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hmbsel][0]_INST_0_i_79_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000808030003000)) 
    \slvi[hmbsel][0]_INST_0_i_8 
       (.I0(hsel326_out),
        .I1(\slvo[4][hconfig][4] [0]),
        .I2(hsel288_in),
        .I3(hsel327_out),
        .I4(\slvi[hmbsel][2]_INST_0_i_9_n_0 ),
        .I5(\slvi[hmbsel][2]_INST_0_i_10_n_0 ),
        .O(\slvi[hmbsel][0]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_80 
       (.I0(\slvo[6][hconfig][4] [11]),
        .I1(\slvo[6][hconfig][4] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[6][hconfig][4] [12]),
        .I4(\slvo[6][hconfig][4] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hmbsel][0]_INST_0_i_80_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_81 
       (.I0(\slvo[6][hconfig][4] [8]),
        .I1(\slvo[6][hconfig][4] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[6][hconfig][4] [9]),
        .I4(\slvo[6][hconfig][4] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hmbsel][0]_INST_0_i_81_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_82 
       (.I0(\slvo[6][hconfig][4] [5]),
        .I1(\slvo[6][hconfig][4] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[6][hconfig][4] [6]),
        .I4(\slvo[6][hconfig][4] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hmbsel][0]_INST_0_i_82_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_83 
       (.I0(\slvo[6][hconfig][4] [14]),
        .I1(\slvo[6][hconfig][4] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[6][hconfig][4] [15]),
        .I4(\slvo[6][hconfig][4] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hmbsel][0]_INST_0_i_83_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_84 
       (.I0(\slvo[6][hconfig][4] [11]),
        .I1(\slvo[6][hconfig][4] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[6][hconfig][4] [12]),
        .I4(\slvo[6][hconfig][4] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hmbsel][0]_INST_0_i_84_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_85 
       (.I0(\slvo[6][hconfig][4] [8]),
        .I1(\slvo[6][hconfig][4] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[6][hconfig][4] [9]),
        .I4(\slvo[6][hconfig][4] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hmbsel][0]_INST_0_i_85_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_86 
       (.I0(\slvo[6][hconfig][4] [5]),
        .I1(\slvo[6][hconfig][4] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[6][hconfig][4] [6]),
        .I4(\slvo[6][hconfig][4] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hmbsel][0]_INST_0_i_86_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_87 
       (.I0(\slvo[4][hconfig][4] [14]),
        .I1(\slvo[4][hconfig][4] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[4][hconfig][4] [15]),
        .I4(\slvo[4][hconfig][4] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hmbsel][0]_INST_0_i_87_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_88 
       (.I0(\slvo[4][hconfig][4] [11]),
        .I1(\slvo[4][hconfig][4] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[4][hconfig][4] [12]),
        .I4(\slvo[4][hconfig][4] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hmbsel][0]_INST_0_i_88_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_89 
       (.I0(\slvo[4][hconfig][4] [8]),
        .I1(\slvo[4][hconfig][4] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[4][hconfig][4] [9]),
        .I4(\slvo[4][hconfig][4] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hmbsel][0]_INST_0_i_89_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \slvi[hmbsel][0]_INST_0_i_9 
       (.I0(hsel2168_in),
        .I1(hsel359_out),
        .I2(hsel330_in),
        .O(hsel1171_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_90 
       (.I0(\slvo[4][hconfig][4] [5]),
        .I1(\slvo[4][hconfig][4] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[4][hconfig][4] [6]),
        .I4(\slvo[4][hconfig][4] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hmbsel][0]_INST_0_i_90_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_91 
       (.I0(\slvo[4][hconfig][4] [14]),
        .I1(\slvo[4][hconfig][4] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[4][hconfig][4] [15]),
        .I4(\slvo[4][hconfig][4] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hmbsel][0]_INST_0_i_91_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_92 
       (.I0(\slvo[4][hconfig][4] [11]),
        .I1(\slvo[4][hconfig][4] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[4][hconfig][4] [12]),
        .I4(\slvo[4][hconfig][4] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hmbsel][0]_INST_0_i_92_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_93 
       (.I0(\slvo[4][hconfig][4] [8]),
        .I1(\slvo[4][hconfig][4] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[4][hconfig][4] [9]),
        .I4(\slvo[4][hconfig][4] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hmbsel][0]_INST_0_i_93_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_94 
       (.I0(\slvo[4][hconfig][4] [5]),
        .I1(\slvo[4][hconfig][4] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[4][hconfig][4] [6]),
        .I4(\slvo[4][hconfig][4] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hmbsel][0]_INST_0_i_94_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_95 
       (.I0(\slvo[3][hconfig][4] [14]),
        .I1(\slvo[3][hconfig][4] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[3][hconfig][4] [15]),
        .I4(\slvo[3][hconfig][4] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hmbsel][0]_INST_0_i_95_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_96 
       (.I0(\slvo[3][hconfig][4] [11]),
        .I1(\slvo[3][hconfig][4] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[3][hconfig][4] [12]),
        .I4(\slvo[3][hconfig][4] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hmbsel][0]_INST_0_i_96_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_97 
       (.I0(\slvo[3][hconfig][4] [8]),
        .I1(\slvo[3][hconfig][4] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[3][hconfig][4] [9]),
        .I4(\slvo[3][hconfig][4] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hmbsel][0]_INST_0_i_97_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_98 
       (.I0(\slvo[3][hconfig][4] [5]),
        .I1(\slvo[3][hconfig][4] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[3][hconfig][4] [6]),
        .I4(\slvo[3][hconfig][4] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hmbsel][0]_INST_0_i_98_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][0]_INST_0_i_99 
       (.I0(\slvo[3][hconfig][4] [14]),
        .I1(\slvo[3][hconfig][4] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[3][hconfig][4] [15]),
        .I4(\slvo[3][hconfig][4] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hmbsel][0]_INST_0_i_99_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF7FFFFFFFFFFFFFF)) 
    \slvi[hmbsel][1]_INST_0 
       (.I0(\slvi[hmbsel][1]_INST_0_i_1_n_0 ),
        .I1(\slvi[hmbsel][1]_INST_0_i_2_n_0 ),
        .I2(\slvi[hmbsel][1]_INST_0_i_3_n_0 ),
        .I3(\slvi[hmbsel][1]_INST_0_i_4_n_0 ),
        .I4(\slvi[hmbsel][1]_INST_0_i_5_n_0 ),
        .I5(\slvi[hmbsel][1]_INST_0_i_6_n_0 ),
        .O(\slvi[hmbsel] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][1]_INST_0_i_1 
       (.I0(\slvo[6][hconfig][5] [1]),
        .I1(\slvi[hmbsel][1]_INST_0_i_7_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000808030003000)) 
    \slvi[hmbsel][1]_INST_0_i_10 
       (.I0(hsel317_out),
        .I1(\slvo[5][hconfig][5] [0]),
        .I2(hsel265_in),
        .I3(hsel320_out),
        .I4(\slvi[hmbsel][2]_INST_0_i_9_n_0 ),
        .I5(\slvi[hmbsel][2]_INST_0_i_10_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_100 
       (.I0(\slvo[3][hconfig][5] [5]),
        .I1(\slvo[3][hconfig][5] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[3][hconfig][5] [6]),
        .I4(\slvo[3][hconfig][5] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hmbsel][1]_INST_0_i_100_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_101 
       (.I0(\slvo[5][hconfig][5] [14]),
        .I1(\slvo[5][hconfig][5] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[5][hconfig][5] [15]),
        .I4(\slvo[5][hconfig][5] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hmbsel][1]_INST_0_i_101_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_102 
       (.I0(\slvo[5][hconfig][5] [11]),
        .I1(\slvo[5][hconfig][5] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[5][hconfig][5] [12]),
        .I4(\slvo[5][hconfig][5] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hmbsel][1]_INST_0_i_102_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_103 
       (.I0(\slvo[5][hconfig][5] [8]),
        .I1(\slvo[5][hconfig][5] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[5][hconfig][5] [9]),
        .I4(\slvo[5][hconfig][5] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hmbsel][1]_INST_0_i_103_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_104 
       (.I0(\slvo[5][hconfig][5] [5]),
        .I1(\slvo[5][hconfig][5] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[5][hconfig][5] [6]),
        .I4(\slvo[5][hconfig][5] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hmbsel][1]_INST_0_i_104_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_105 
       (.I0(\slvo[5][hconfig][5] [14]),
        .I1(\slvo[5][hconfig][5] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[5][hconfig][5] [15]),
        .I4(\slvo[5][hconfig][5] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hmbsel][1]_INST_0_i_105_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_106 
       (.I0(\slvo[5][hconfig][5] [11]),
        .I1(\slvo[5][hconfig][5] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[5][hconfig][5] [12]),
        .I4(\slvo[5][hconfig][5] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hmbsel][1]_INST_0_i_106_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_107 
       (.I0(\slvo[5][hconfig][5] [8]),
        .I1(\slvo[5][hconfig][5] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[5][hconfig][5] [9]),
        .I4(\slvo[5][hconfig][5] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hmbsel][1]_INST_0_i_107_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_108 
       (.I0(\slvo[5][hconfig][5] [5]),
        .I1(\slvo[5][hconfig][5] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[5][hconfig][5] [6]),
        .I4(\slvo[5][hconfig][5] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hmbsel][1]_INST_0_i_108_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_109 
       (.I0(\slvo[7][hconfig][5] [14]),
        .I1(\slvo[7][hconfig][5] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[7][hconfig][5] [15]),
        .I4(\slvo[7][hconfig][5] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hmbsel][1]_INST_0_i_109_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000808030003000)) 
    \slvi[hmbsel][1]_INST_0_i_11 
       (.I0(hsel31_out),
        .I1(\slvo[7][hconfig][5] [0]),
        .I2(hsel224_in),
        .I3(hsel34_out),
        .I4(\slvi[hmbsel][2]_INST_0_i_9_n_0 ),
        .I5(\slvi[hmbsel][2]_INST_0_i_10_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_110 
       (.I0(\slvo[7][hconfig][5] [11]),
        .I1(\slvo[7][hconfig][5] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[7][hconfig][5] [12]),
        .I4(\slvo[7][hconfig][5] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hmbsel][1]_INST_0_i_110_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_111 
       (.I0(\slvo[7][hconfig][5] [8]),
        .I1(\slvo[7][hconfig][5] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[7][hconfig][5] [9]),
        .I4(\slvo[7][hconfig][5] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hmbsel][1]_INST_0_i_111_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_112 
       (.I0(\slvo[7][hconfig][5] [5]),
        .I1(\slvo[7][hconfig][5] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[7][hconfig][5] [6]),
        .I4(\slvo[7][hconfig][5] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hmbsel][1]_INST_0_i_112_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_113 
       (.I0(\slvo[7][hconfig][5] [14]),
        .I1(\slvo[7][hconfig][5] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[7][hconfig][5] [15]),
        .I4(\slvo[7][hconfig][5] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hmbsel][1]_INST_0_i_113_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_114 
       (.I0(\slvo[7][hconfig][5] [11]),
        .I1(\slvo[7][hconfig][5] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[7][hconfig][5] [12]),
        .I4(\slvo[7][hconfig][5] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hmbsel][1]_INST_0_i_114_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_115 
       (.I0(\slvo[7][hconfig][5] [8]),
        .I1(\slvo[7][hconfig][5] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[7][hconfig][5] [9]),
        .I4(\slvo[7][hconfig][5] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hmbsel][1]_INST_0_i_115_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_116 
       (.I0(\slvo[7][hconfig][5] [5]),
        .I1(\slvo[7][hconfig][5] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[7][hconfig][5] [6]),
        .I4(\slvo[7][hconfig][5] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hmbsel][1]_INST_0_i_116_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][1]_INST_0_i_12 
       (.CI(slvi),
        .CO({hsel39_out,\slvi[hmbsel][1]_INST_0_i_12_n_1 ,\slvi[hmbsel][1]_INST_0_i_12_n_2 ,\slvi[hmbsel][1]_INST_0_i_12_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][1]_INST_0_i_27_n_0 ,\slvi[hmbsel][1]_INST_0_i_28_n_0 ,\slvi[hmbsel][1]_INST_0_i_29_n_0 ,\slvi[hmbsel][1]_INST_0_i_30_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][1]_INST_0_i_13 
       (.I0(\slvi[hmbsel][1]_INST_0_i_31_n_0 ),
        .I1(\slvi[hmbsel][1]_INST_0_i_32_n_0 ),
        .O(hsel245_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][1]_INST_0_i_14 
       (.CI(slvi),
        .CO({hsel312_out,\slvi[hmbsel][1]_INST_0_i_14_n_1 ,\slvi[hmbsel][1]_INST_0_i_14_n_2 ,\slvi[hmbsel][1]_INST_0_i_14_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][1]_INST_0_i_33_n_0 ,\slvi[hmbsel][1]_INST_0_i_34_n_0 ,\slvi[hmbsel][1]_INST_0_i_35_n_0 ,\slvi[hmbsel][1]_INST_0_i_36_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][1]_INST_0_i_15 
       (.CI(slvi),
        .CO({hsel325_out,\slvi[hmbsel][1]_INST_0_i_15_n_1 ,\slvi[hmbsel][1]_INST_0_i_15_n_2 ,\slvi[hmbsel][1]_INST_0_i_15_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][1]_INST_0_i_37_n_0 ,\slvi[hmbsel][1]_INST_0_i_38_n_0 ,\slvi[hmbsel][1]_INST_0_i_39_n_0 ,\slvi[hmbsel][1]_INST_0_i_40_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][1]_INST_0_i_16 
       (.I0(\slvi[hmbsel][1]_INST_0_i_41_n_0 ),
        .I1(\slvi[hmbsel][1]_INST_0_i_42_n_0 ),
        .O(hsel285_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][1]_INST_0_i_17 
       (.CI(slvi),
        .CO({hsel328_out,\slvi[hmbsel][1]_INST_0_i_17_n_1 ,\slvi[hmbsel][1]_INST_0_i_17_n_2 ,\slvi[hmbsel][1]_INST_0_i_17_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][1]_INST_0_i_43_n_0 ,\slvi[hmbsel][1]_INST_0_i_44_n_0 ,\slvi[hmbsel][1]_INST_0_i_45_n_0 ,\slvi[hmbsel][1]_INST_0_i_46_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][1]_INST_0_i_18 
       (.CI(slvi),
        .CO({hsel333_out,\slvi[hmbsel][1]_INST_0_i_18_n_1 ,\slvi[hmbsel][1]_INST_0_i_18_n_2 ,\slvi[hmbsel][1]_INST_0_i_18_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][1]_INST_0_i_47_n_0 ,\slvi[hmbsel][1]_INST_0_i_48_n_0 ,\slvi[hmbsel][1]_INST_0_i_49_n_0 ,\slvi[hmbsel][1]_INST_0_i_50_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][1]_INST_0_i_19 
       (.I0(\slvi[hmbsel][1]_INST_0_i_51_n_0 ),
        .I1(\slvi[hmbsel][1]_INST_0_i_52_n_0 ),
        .O(hsel2105_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][1]_INST_0_i_2 
       (.I0(\slvo[4][hconfig][5] [1]),
        .I1(\slvi[hmbsel][1]_INST_0_i_8_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][1]_INST_0_i_20 
       (.CI(slvi),
        .CO({hsel336_out,\slvi[hmbsel][1]_INST_0_i_20_n_1 ,\slvi[hmbsel][1]_INST_0_i_20_n_2 ,\slvi[hmbsel][1]_INST_0_i_20_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][1]_INST_0_i_53_n_0 ,\slvi[hmbsel][1]_INST_0_i_54_n_0 ,\slvi[hmbsel][1]_INST_0_i_55_n_0 ,\slvi[hmbsel][1]_INST_0_i_56_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][1]_INST_0_i_21 
       (.CI(slvi),
        .CO({hsel317_out,\slvi[hmbsel][1]_INST_0_i_21_n_1 ,\slvi[hmbsel][1]_INST_0_i_21_n_2 ,\slvi[hmbsel][1]_INST_0_i_21_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][1]_INST_0_i_57_n_0 ,\slvi[hmbsel][1]_INST_0_i_58_n_0 ,\slvi[hmbsel][1]_INST_0_i_59_n_0 ,\slvi[hmbsel][1]_INST_0_i_60_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][1]_INST_0_i_22 
       (.I0(\slvi[hmbsel][1]_INST_0_i_61_n_0 ),
        .I1(\slvi[hmbsel][1]_INST_0_i_62_n_0 ),
        .O(hsel265_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][1]_INST_0_i_23 
       (.CI(slvi),
        .CO({hsel320_out,\slvi[hmbsel][1]_INST_0_i_23_n_1 ,\slvi[hmbsel][1]_INST_0_i_23_n_2 ,\slvi[hmbsel][1]_INST_0_i_23_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][1]_INST_0_i_63_n_0 ,\slvi[hmbsel][1]_INST_0_i_64_n_0 ,\slvi[hmbsel][1]_INST_0_i_65_n_0 ,\slvi[hmbsel][1]_INST_0_i_66_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][1]_INST_0_i_24 
       (.CI(slvi),
        .CO({hsel31_out,\slvi[hmbsel][1]_INST_0_i_24_n_1 ,\slvi[hmbsel][1]_INST_0_i_24_n_2 ,\slvi[hmbsel][1]_INST_0_i_24_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][1]_INST_0_i_67_n_0 ,\slvi[hmbsel][1]_INST_0_i_68_n_0 ,\slvi[hmbsel][1]_INST_0_i_69_n_0 ,\slvi[hmbsel][1]_INST_0_i_70_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][1]_INST_0_i_25 
       (.I0(\slvi[hmbsel][1]_INST_0_i_71_n_0 ),
        .I1(\slvi[hmbsel][1]_INST_0_i_72_n_0 ),
        .O(hsel224_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][1]_INST_0_i_26 
       (.CI(slvi),
        .CO({hsel34_out,\slvi[hmbsel][1]_INST_0_i_26_n_1 ,\slvi[hmbsel][1]_INST_0_i_26_n_2 ,\slvi[hmbsel][1]_INST_0_i_26_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][1]_INST_0_i_73_n_0 ,\slvi[hmbsel][1]_INST_0_i_74_n_0 ,\slvi[hmbsel][1]_INST_0_i_75_n_0 ,\slvi[hmbsel][1]_INST_0_i_76_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_27 
       (.I0(\slvo[6][hconfig][5] [13]),
        .I1(\slvo[6][hconfig][5] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hmbsel][1]_INST_0_i_77_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_28 
       (.I0(\slvo[6][hconfig][5] [10]),
        .I1(\slvo[6][hconfig][5] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hmbsel][1]_INST_0_i_78_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_29 
       (.I0(\slvo[6][hconfig][5] [7]),
        .I1(\slvo[6][hconfig][5] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hmbsel][1]_INST_0_i_79_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFD5D5555FFFFFFFF)) 
    \slvi[hmbsel][1]_INST_0_i_3 
       (.I0(\slvi[hsel][1]_INST_0_i_3_n_0 ),
        .I1(hsel1173_out),
        .I2(\slvo[0][hconfig][5] [0]),
        .I3(hsel1166_out),
        .I4(\slvo[0][hconfig][5] [1]),
        .I5(\slvi[hsel][2]_INST_0_i_2_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_30 
       (.I0(\slvo[6][hconfig][5] [4]),
        .I1(\slvo[6][hconfig][5] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hmbsel][1]_INST_0_i_80_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][1]_INST_0_i_31 
       (.I0(\slvo[6][hconfig][5] [9]),
        .I1(\slvo[6][hconfig][5] [7]),
        .I2(\slvo[6][hconfig][5] [8]),
        .I3(\slvo[6][hconfig][5] [4]),
        .I4(\slvo[6][hconfig][5] [5]),
        .I5(\slvo[6][hconfig][5] [6]),
        .O(\slvi[hmbsel][1]_INST_0_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][1]_INST_0_i_32 
       (.I0(\slvo[6][hconfig][5] [14]),
        .I1(\slvo[6][hconfig][5] [13]),
        .I2(\slvo[6][hconfig][5] [15]),
        .I3(\slvo[6][hconfig][5] [10]),
        .I4(\slvo[6][hconfig][5] [11]),
        .I5(\slvo[6][hconfig][5] [12]),
        .O(\slvi[hmbsel][1]_INST_0_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_33 
       (.I0(\slvo[6][hconfig][5] [13]),
        .I1(\slvo[6][hconfig][5] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hmbsel][1]_INST_0_i_81_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_34 
       (.I0(\slvo[6][hconfig][5] [10]),
        .I1(\slvo[6][hconfig][5] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hmbsel][1]_INST_0_i_82_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_35 
       (.I0(\slvo[6][hconfig][5] [7]),
        .I1(\slvo[6][hconfig][5] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hmbsel][1]_INST_0_i_83_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_36 
       (.I0(\slvo[6][hconfig][5] [4]),
        .I1(\slvo[6][hconfig][5] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hmbsel][1]_INST_0_i_84_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_37 
       (.I0(\slvo[4][hconfig][5] [13]),
        .I1(\slvo[4][hconfig][5] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hmbsel][1]_INST_0_i_85_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_38 
       (.I0(\slvo[4][hconfig][5] [10]),
        .I1(\slvo[4][hconfig][5] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hmbsel][1]_INST_0_i_86_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_39 
       (.I0(\slvo[4][hconfig][5] [7]),
        .I1(\slvo[4][hconfig][5] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hmbsel][1]_INST_0_i_87_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][1]_INST_0_i_4 
       (.I0(\slvo[3][hconfig][5] [1]),
        .I1(\slvi[hmbsel][1]_INST_0_i_9_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_40 
       (.I0(\slvo[4][hconfig][5] [4]),
        .I1(\slvo[4][hconfig][5] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hmbsel][1]_INST_0_i_88_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][1]_INST_0_i_41 
       (.I0(\slvo[4][hconfig][5] [9]),
        .I1(\slvo[4][hconfig][5] [7]),
        .I2(\slvo[4][hconfig][5] [8]),
        .I3(\slvo[4][hconfig][5] [4]),
        .I4(\slvo[4][hconfig][5] [5]),
        .I5(\slvo[4][hconfig][5] [6]),
        .O(\slvi[hmbsel][1]_INST_0_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][1]_INST_0_i_42 
       (.I0(\slvo[4][hconfig][5] [14]),
        .I1(\slvo[4][hconfig][5] [13]),
        .I2(\slvo[4][hconfig][5] [15]),
        .I3(\slvo[4][hconfig][5] [10]),
        .I4(\slvo[4][hconfig][5] [11]),
        .I5(\slvo[4][hconfig][5] [12]),
        .O(\slvi[hmbsel][1]_INST_0_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_43 
       (.I0(\slvo[4][hconfig][5] [13]),
        .I1(\slvo[4][hconfig][5] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hmbsel][1]_INST_0_i_89_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_44 
       (.I0(\slvo[4][hconfig][5] [10]),
        .I1(\slvo[4][hconfig][5] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hmbsel][1]_INST_0_i_90_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_45 
       (.I0(\slvo[4][hconfig][5] [7]),
        .I1(\slvo[4][hconfig][5] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hmbsel][1]_INST_0_i_91_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_46 
       (.I0(\slvo[4][hconfig][5] [4]),
        .I1(\slvo[4][hconfig][5] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hmbsel][1]_INST_0_i_92_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_47 
       (.I0(\slvo[3][hconfig][5] [13]),
        .I1(\slvo[3][hconfig][5] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hmbsel][1]_INST_0_i_93_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_48 
       (.I0(\slvo[3][hconfig][5] [10]),
        .I1(\slvo[3][hconfig][5] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hmbsel][1]_INST_0_i_94_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_49 
       (.I0(\slvo[3][hconfig][5] [7]),
        .I1(\slvo[3][hconfig][5] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hmbsel][1]_INST_0_i_95_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][1]_INST_0_i_5 
       (.I0(\slvo[5][hconfig][5] [1]),
        .I1(\slvi[hmbsel][1]_INST_0_i_10_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_50 
       (.I0(\slvo[3][hconfig][5] [4]),
        .I1(\slvo[3][hconfig][5] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hmbsel][1]_INST_0_i_96_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][1]_INST_0_i_51 
       (.I0(\slvo[3][hconfig][5] [9]),
        .I1(\slvo[3][hconfig][5] [7]),
        .I2(\slvo[3][hconfig][5] [8]),
        .I3(\slvo[3][hconfig][5] [4]),
        .I4(\slvo[3][hconfig][5] [5]),
        .I5(\slvo[3][hconfig][5] [6]),
        .O(\slvi[hmbsel][1]_INST_0_i_51_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][1]_INST_0_i_52 
       (.I0(\slvo[3][hconfig][5] [14]),
        .I1(\slvo[3][hconfig][5] [13]),
        .I2(\slvo[3][hconfig][5] [15]),
        .I3(\slvo[3][hconfig][5] [10]),
        .I4(\slvo[3][hconfig][5] [11]),
        .I5(\slvo[3][hconfig][5] [12]),
        .O(\slvi[hmbsel][1]_INST_0_i_52_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_53 
       (.I0(\slvo[3][hconfig][5] [13]),
        .I1(\slvo[3][hconfig][5] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hmbsel][1]_INST_0_i_97_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_53_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_54 
       (.I0(\slvo[3][hconfig][5] [10]),
        .I1(\slvo[3][hconfig][5] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hmbsel][1]_INST_0_i_98_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_54_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_55 
       (.I0(\slvo[3][hconfig][5] [7]),
        .I1(\slvo[3][hconfig][5] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hmbsel][1]_INST_0_i_99_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_55_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_56 
       (.I0(\slvo[3][hconfig][5] [4]),
        .I1(\slvo[3][hconfig][5] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hmbsel][1]_INST_0_i_100_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_56_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_57 
       (.I0(\slvo[5][hconfig][5] [13]),
        .I1(\slvo[5][hconfig][5] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hmbsel][1]_INST_0_i_101_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_57_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_58 
       (.I0(\slvo[5][hconfig][5] [10]),
        .I1(\slvo[5][hconfig][5] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hmbsel][1]_INST_0_i_102_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_58_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_59 
       (.I0(\slvo[5][hconfig][5] [7]),
        .I1(\slvo[5][hconfig][5] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hmbsel][1]_INST_0_i_103_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_59_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][1]_INST_0_i_6 
       (.I0(\slvo[7][hconfig][5] [1]),
        .I1(\slvi[hmbsel][1]_INST_0_i_11_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_60 
       (.I0(\slvo[5][hconfig][5] [4]),
        .I1(\slvo[5][hconfig][5] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hmbsel][1]_INST_0_i_104_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_60_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][1]_INST_0_i_61 
       (.I0(\slvo[5][hconfig][5] [9]),
        .I1(\slvo[5][hconfig][5] [7]),
        .I2(\slvo[5][hconfig][5] [8]),
        .I3(\slvo[5][hconfig][5] [4]),
        .I4(\slvo[5][hconfig][5] [5]),
        .I5(\slvo[5][hconfig][5] [6]),
        .O(\slvi[hmbsel][1]_INST_0_i_61_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][1]_INST_0_i_62 
       (.I0(\slvo[5][hconfig][5] [14]),
        .I1(\slvo[5][hconfig][5] [13]),
        .I2(\slvo[5][hconfig][5] [15]),
        .I3(\slvo[5][hconfig][5] [10]),
        .I4(\slvo[5][hconfig][5] [11]),
        .I5(\slvo[5][hconfig][5] [12]),
        .O(\slvi[hmbsel][1]_INST_0_i_62_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_63 
       (.I0(\slvo[5][hconfig][5] [13]),
        .I1(\slvo[5][hconfig][5] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hmbsel][1]_INST_0_i_105_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_63_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_64 
       (.I0(\slvo[5][hconfig][5] [10]),
        .I1(\slvo[5][hconfig][5] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hmbsel][1]_INST_0_i_106_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_64_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_65 
       (.I0(\slvo[5][hconfig][5] [7]),
        .I1(\slvo[5][hconfig][5] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hmbsel][1]_INST_0_i_107_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_65_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_66 
       (.I0(\slvo[5][hconfig][5] [4]),
        .I1(\slvo[5][hconfig][5] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hmbsel][1]_INST_0_i_108_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_66_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_67 
       (.I0(\slvo[7][hconfig][5] [13]),
        .I1(\slvo[7][hconfig][5] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hmbsel][1]_INST_0_i_109_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_67_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_68 
       (.I0(\slvo[7][hconfig][5] [10]),
        .I1(\slvo[7][hconfig][5] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hmbsel][1]_INST_0_i_110_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_68_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_69 
       (.I0(\slvo[7][hconfig][5] [7]),
        .I1(\slvo[7][hconfig][5] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hmbsel][1]_INST_0_i_111_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_69_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000808030003000)) 
    \slvi[hmbsel][1]_INST_0_i_7 
       (.I0(hsel39_out),
        .I1(\slvo[6][hconfig][5] [0]),
        .I2(hsel245_in),
        .I3(hsel312_out),
        .I4(\slvi[hmbsel][2]_INST_0_i_9_n_0 ),
        .I5(\slvi[hmbsel][2]_INST_0_i_10_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_70 
       (.I0(\slvo[7][hconfig][5] [4]),
        .I1(\slvo[7][hconfig][5] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hmbsel][1]_INST_0_i_112_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_70_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][1]_INST_0_i_71 
       (.I0(\slvo[7][hconfig][5] [9]),
        .I1(\slvo[7][hconfig][5] [7]),
        .I2(\slvo[7][hconfig][5] [8]),
        .I3(\slvo[7][hconfig][5] [4]),
        .I4(\slvo[7][hconfig][5] [5]),
        .I5(\slvo[7][hconfig][5] [6]),
        .O(\slvi[hmbsel][1]_INST_0_i_71_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][1]_INST_0_i_72 
       (.I0(\slvo[7][hconfig][5] [14]),
        .I1(\slvo[7][hconfig][5] [13]),
        .I2(\slvo[7][hconfig][5] [15]),
        .I3(\slvo[7][hconfig][5] [10]),
        .I4(\slvo[7][hconfig][5] [11]),
        .I5(\slvo[7][hconfig][5] [12]),
        .O(\slvi[hmbsel][1]_INST_0_i_72_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_73 
       (.I0(\slvo[7][hconfig][5] [13]),
        .I1(\slvo[7][hconfig][5] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hmbsel][1]_INST_0_i_113_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_73_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_74 
       (.I0(\slvo[7][hconfig][5] [10]),
        .I1(\slvo[7][hconfig][5] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hmbsel][1]_INST_0_i_114_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_74_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_75 
       (.I0(\slvo[7][hconfig][5] [7]),
        .I1(\slvo[7][hconfig][5] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hmbsel][1]_INST_0_i_115_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_75_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][1]_INST_0_i_76 
       (.I0(\slvo[7][hconfig][5] [4]),
        .I1(\slvo[7][hconfig][5] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hmbsel][1]_INST_0_i_116_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_76_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_77 
       (.I0(\slvo[6][hconfig][5] [14]),
        .I1(\slvo[6][hconfig][5] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[6][hconfig][5] [15]),
        .I4(\slvo[6][hconfig][5] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hmbsel][1]_INST_0_i_77_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_78 
       (.I0(\slvo[6][hconfig][5] [11]),
        .I1(\slvo[6][hconfig][5] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[6][hconfig][5] [12]),
        .I4(\slvo[6][hconfig][5] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hmbsel][1]_INST_0_i_78_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_79 
       (.I0(\slvo[6][hconfig][5] [8]),
        .I1(\slvo[6][hconfig][5] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[6][hconfig][5] [9]),
        .I4(\slvo[6][hconfig][5] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hmbsel][1]_INST_0_i_79_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000808030003000)) 
    \slvi[hmbsel][1]_INST_0_i_8 
       (.I0(hsel325_out),
        .I1(\slvo[4][hconfig][5] [0]),
        .I2(hsel285_in),
        .I3(hsel328_out),
        .I4(\slvi[hmbsel][2]_INST_0_i_9_n_0 ),
        .I5(\slvi[hmbsel][2]_INST_0_i_10_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_80 
       (.I0(\slvo[6][hconfig][5] [5]),
        .I1(\slvo[6][hconfig][5] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[6][hconfig][5] [6]),
        .I4(\slvo[6][hconfig][5] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hmbsel][1]_INST_0_i_80_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_81 
       (.I0(\slvo[6][hconfig][5] [14]),
        .I1(\slvo[6][hconfig][5] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[6][hconfig][5] [15]),
        .I4(\slvo[6][hconfig][5] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hmbsel][1]_INST_0_i_81_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_82 
       (.I0(\slvo[6][hconfig][5] [11]),
        .I1(\slvo[6][hconfig][5] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[6][hconfig][5] [12]),
        .I4(\slvo[6][hconfig][5] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hmbsel][1]_INST_0_i_82_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_83 
       (.I0(\slvo[6][hconfig][5] [8]),
        .I1(\slvo[6][hconfig][5] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[6][hconfig][5] [9]),
        .I4(\slvo[6][hconfig][5] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hmbsel][1]_INST_0_i_83_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_84 
       (.I0(\slvo[6][hconfig][5] [5]),
        .I1(\slvo[6][hconfig][5] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[6][hconfig][5] [6]),
        .I4(\slvo[6][hconfig][5] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hmbsel][1]_INST_0_i_84_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_85 
       (.I0(\slvo[4][hconfig][5] [14]),
        .I1(\slvo[4][hconfig][5] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[4][hconfig][5] [15]),
        .I4(\slvo[4][hconfig][5] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hmbsel][1]_INST_0_i_85_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_86 
       (.I0(\slvo[4][hconfig][5] [11]),
        .I1(\slvo[4][hconfig][5] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[4][hconfig][5] [12]),
        .I4(\slvo[4][hconfig][5] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hmbsel][1]_INST_0_i_86_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_87 
       (.I0(\slvo[4][hconfig][5] [8]),
        .I1(\slvo[4][hconfig][5] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[4][hconfig][5] [9]),
        .I4(\slvo[4][hconfig][5] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hmbsel][1]_INST_0_i_87_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_88 
       (.I0(\slvo[4][hconfig][5] [5]),
        .I1(\slvo[4][hconfig][5] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[4][hconfig][5] [6]),
        .I4(\slvo[4][hconfig][5] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hmbsel][1]_INST_0_i_88_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_89 
       (.I0(\slvo[4][hconfig][5] [14]),
        .I1(\slvo[4][hconfig][5] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[4][hconfig][5] [15]),
        .I4(\slvo[4][hconfig][5] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hmbsel][1]_INST_0_i_89_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000808030003000)) 
    \slvi[hmbsel][1]_INST_0_i_9 
       (.I0(hsel333_out),
        .I1(\slvo[3][hconfig][5] [0]),
        .I2(hsel2105_in),
        .I3(hsel336_out),
        .I4(\slvi[hmbsel][2]_INST_0_i_9_n_0 ),
        .I5(\slvi[hmbsel][2]_INST_0_i_10_n_0 ),
        .O(\slvi[hmbsel][1]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_90 
       (.I0(\slvo[4][hconfig][5] [11]),
        .I1(\slvo[4][hconfig][5] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[4][hconfig][5] [12]),
        .I4(\slvo[4][hconfig][5] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hmbsel][1]_INST_0_i_90_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_91 
       (.I0(\slvo[4][hconfig][5] [8]),
        .I1(\slvo[4][hconfig][5] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[4][hconfig][5] [9]),
        .I4(\slvo[4][hconfig][5] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hmbsel][1]_INST_0_i_91_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_92 
       (.I0(\slvo[4][hconfig][5] [5]),
        .I1(\slvo[4][hconfig][5] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[4][hconfig][5] [6]),
        .I4(\slvo[4][hconfig][5] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hmbsel][1]_INST_0_i_92_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_93 
       (.I0(\slvo[3][hconfig][5] [14]),
        .I1(\slvo[3][hconfig][5] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[3][hconfig][5] [15]),
        .I4(\slvo[3][hconfig][5] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hmbsel][1]_INST_0_i_93_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_94 
       (.I0(\slvo[3][hconfig][5] [11]),
        .I1(\slvo[3][hconfig][5] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[3][hconfig][5] [12]),
        .I4(\slvo[3][hconfig][5] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hmbsel][1]_INST_0_i_94_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_95 
       (.I0(\slvo[3][hconfig][5] [8]),
        .I1(\slvo[3][hconfig][5] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[3][hconfig][5] [9]),
        .I4(\slvo[3][hconfig][5] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hmbsel][1]_INST_0_i_95_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_96 
       (.I0(\slvo[3][hconfig][5] [5]),
        .I1(\slvo[3][hconfig][5] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[3][hconfig][5] [6]),
        .I4(\slvo[3][hconfig][5] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hmbsel][1]_INST_0_i_96_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_97 
       (.I0(\slvo[3][hconfig][5] [14]),
        .I1(\slvo[3][hconfig][5] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[3][hconfig][5] [15]),
        .I4(\slvo[3][hconfig][5] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hmbsel][1]_INST_0_i_97_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_98 
       (.I0(\slvo[3][hconfig][5] [11]),
        .I1(\slvo[3][hconfig][5] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[3][hconfig][5] [12]),
        .I4(\slvo[3][hconfig][5] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hmbsel][1]_INST_0_i_98_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][1]_INST_0_i_99 
       (.I0(\slvo[3][hconfig][5] [8]),
        .I1(\slvo[3][hconfig][5] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[3][hconfig][5] [9]),
        .I4(\slvo[3][hconfig][5] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hmbsel][1]_INST_0_i_99_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \slvi[hmbsel][2]_INST_0 
       (.I0(\slvo[7][hconfig][6] [1]),
        .I1(\slvi[hmbsel][2]_INST_0_i_1_n_0 ),
        .I2(\slvi[hmbsel][2]_INST_0_i_2_n_0 ),
        .I3(\slvi[hmbsel][2]_INST_0_i_3_n_0 ),
        .I4(\slvi[hmbsel][2]_INST_0_i_4_n_0 ),
        .I5(\slvi[hmbsel][2]_INST_0_i_5_n_0 ),
        .O(\slvi[hmbsel] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000808030003000)) 
    \slvi[hmbsel][2]_INST_0_i_1 
       (.I0(hsel30_out),
        .I1(\slvo[7][hconfig][6] [0]),
        .I2(hsel221_in),
        .I3(hsel35_out),
        .I4(\slvi[hmbsel][2]_INST_0_i_9_n_0 ),
        .I5(\slvi[hmbsel][2]_INST_0_i_10_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \slvi[hmbsel][2]_INST_0_i_10 
       (.I0(\slvi[haddr] [29]),
        .I1(\slvi[haddr] [31]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvi[haddr] [28]),
        .I4(\slvi[haddr] [26]),
        .I5(\slvi[haddr] [27]),
        .O(\slvi[hmbsel][2]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000808030003000)) 
    \slvi[hmbsel][2]_INST_0_i_11 
       (.I0(hsel38_out),
        .I1(\slvo[6][hconfig][6] [0]),
        .I2(hsel242_in),
        .I3(hsel313_out),
        .I4(\slvi[hmbsel][2]_INST_0_i_9_n_0 ),
        .I5(\slvi[hmbsel][2]_INST_0_i_10_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000808030003000)) 
    \slvi[hmbsel][2]_INST_0_i_12 
       (.I0(hsel324_out),
        .I1(\slvo[4][hconfig][6] [0]),
        .I2(hsel282_in),
        .I3(hsel329_out),
        .I4(\slvi[hmbsel][2]_INST_0_i_9_n_0 ),
        .I5(\slvi[hmbsel][2]_INST_0_i_10_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8F00800080008000)) 
    \slvi[hmbsel][2]_INST_0_i_13 
       (.I0(hsel356_out),
        .I1(hsel219_in),
        .I2(\slvo[0][hconfig][6] [0]),
        .I3(hsel2162_in),
        .I4(hsel361_out),
        .I5(hsel330_in),
        .O(\slvi[hmbsel][2]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8F00800080008000)) 
    \slvi[hmbsel][2]_INST_0_i_14 
       (.I0(hsel348_out),
        .I1(hsel219_in),
        .I2(\slvo[1][hconfig][6] [0]),
        .I3(hsel2142_in),
        .I4(hsel353_out),
        .I5(hsel330_in),
        .O(\slvi[hmbsel][2]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000808030003000)) 
    \slvi[hmbsel][2]_INST_0_i_15 
       (.I0(hsel316_out),
        .I1(\slvo[5][hconfig][6] [0]),
        .I2(hsel262_in),
        .I3(hsel321_out),
        .I4(\slvi[hmbsel][2]_INST_0_i_9_n_0 ),
        .I5(\slvi[hmbsel][2]_INST_0_i_10_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_16 
       (.I0(\slvo[7][hconfig][6] [13]),
        .I1(\slvo[7][hconfig][6] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hmbsel][2]_INST_0_i_35_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_17 
       (.I0(\slvo[7][hconfig][6] [10]),
        .I1(\slvo[7][hconfig][6] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hmbsel][2]_INST_0_i_36_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_18 
       (.I0(\slvo[7][hconfig][6] [7]),
        .I1(\slvo[7][hconfig][6] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hmbsel][2]_INST_0_i_37_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_19 
       (.I0(\slvo[7][hconfig][6] [4]),
        .I1(\slvo[7][hconfig][6] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hmbsel][2]_INST_0_i_38_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \slvi[hmbsel][2]_INST_0_i_2 
       (.I0(\slvi[hmbsel][2]_INST_0_i_11_n_0 ),
        .I1(\slvo[6][hconfig][6] [1]),
        .O(\slvi[hmbsel][2]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][2]_INST_0_i_20 
       (.I0(\slvo[7][hconfig][6] [9]),
        .I1(\slvo[7][hconfig][6] [7]),
        .I2(\slvo[7][hconfig][6] [8]),
        .I3(\slvo[7][hconfig][6] [4]),
        .I4(\slvo[7][hconfig][6] [5]),
        .I5(\slvo[7][hconfig][6] [6]),
        .O(\slvi[hmbsel][2]_INST_0_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][2]_INST_0_i_21 
       (.I0(\slvo[7][hconfig][6] [14]),
        .I1(\slvo[7][hconfig][6] [13]),
        .I2(\slvo[7][hconfig][6] [15]),
        .I3(\slvo[7][hconfig][6] [10]),
        .I4(\slvo[7][hconfig][6] [11]),
        .I5(\slvo[7][hconfig][6] [12]),
        .O(\slvi[hmbsel][2]_INST_0_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_22 
       (.I0(\slvo[7][hconfig][6] [13]),
        .I1(\slvo[7][hconfig][6] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hmbsel][2]_INST_0_i_39_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_23 
       (.I0(\slvo[7][hconfig][6] [10]),
        .I1(\slvo[7][hconfig][6] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hmbsel][2]_INST_0_i_40_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_24 
       (.I0(\slvo[7][hconfig][6] [7]),
        .I1(\slvo[7][hconfig][6] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hmbsel][2]_INST_0_i_41_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_25 
       (.I0(\slvo[7][hconfig][6] [4]),
        .I1(\slvo[7][hconfig][6] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hmbsel][2]_INST_0_i_42_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][2]_INST_0_i_26 
       (.CI(slvi),
        .CO({hsel38_out,\slvi[hmbsel][2]_INST_0_i_26_n_1 ,\slvi[hmbsel][2]_INST_0_i_26_n_2 ,\slvi[hmbsel][2]_INST_0_i_26_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][2]_INST_0_i_43_n_0 ,\slvi[hmbsel][2]_INST_0_i_44_n_0 ,\slvi[hmbsel][2]_INST_0_i_45_n_0 ,\slvi[hmbsel][2]_INST_0_i_46_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][2]_INST_0_i_27 
       (.I0(\slvi[hmbsel][2]_INST_0_i_47_n_0 ),
        .I1(\slvi[hmbsel][2]_INST_0_i_48_n_0 ),
        .O(hsel242_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][2]_INST_0_i_28 
       (.CI(slvi),
        .CO({hsel313_out,\slvi[hmbsel][2]_INST_0_i_28_n_1 ,\slvi[hmbsel][2]_INST_0_i_28_n_2 ,\slvi[hmbsel][2]_INST_0_i_28_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][2]_INST_0_i_49_n_0 ,\slvi[hmbsel][2]_INST_0_i_50_n_0 ,\slvi[hmbsel][2]_INST_0_i_51_n_0 ,\slvi[hmbsel][2]_INST_0_i_52_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][2]_INST_0_i_29 
       (.CI(slvi),
        .CO({hsel324_out,\slvi[hmbsel][2]_INST_0_i_29_n_1 ,\slvi[hmbsel][2]_INST_0_i_29_n_2 ,\slvi[hmbsel][2]_INST_0_i_29_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][2]_INST_0_i_53_n_0 ,\slvi[hmbsel][2]_INST_0_i_54_n_0 ,\slvi[hmbsel][2]_INST_0_i_55_n_0 ,\slvi[hmbsel][2]_INST_0_i_56_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \slvi[hmbsel][2]_INST_0_i_3 
       (.I0(\slvi[hmbsel][2]_INST_0_i_12_n_0 ),
        .I1(\slvo[4][hconfig][6] [1]),
        .O(\slvi[hmbsel][2]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][2]_INST_0_i_30 
       (.I0(\slvi[hmbsel][2]_INST_0_i_57_n_0 ),
        .I1(\slvi[hmbsel][2]_INST_0_i_58_n_0 ),
        .O(hsel282_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][2]_INST_0_i_31 
       (.CI(slvi),
        .CO({hsel329_out,\slvi[hmbsel][2]_INST_0_i_31_n_1 ,\slvi[hmbsel][2]_INST_0_i_31_n_2 ,\slvi[hmbsel][2]_INST_0_i_31_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][2]_INST_0_i_59_n_0 ,\slvi[hmbsel][2]_INST_0_i_60_n_0 ,\slvi[hmbsel][2]_INST_0_i_61_n_0 ,\slvi[hmbsel][2]_INST_0_i_62_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][2]_INST_0_i_32 
       (.CI(slvi),
        .CO({hsel316_out,\slvi[hmbsel][2]_INST_0_i_32_n_1 ,\slvi[hmbsel][2]_INST_0_i_32_n_2 ,\slvi[hmbsel][2]_INST_0_i_32_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][2]_INST_0_i_63_n_0 ,\slvi[hmbsel][2]_INST_0_i_64_n_0 ,\slvi[hmbsel][2]_INST_0_i_65_n_0 ,\slvi[hmbsel][2]_INST_0_i_66_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][2]_INST_0_i_33 
       (.I0(\slvi[hmbsel][2]_INST_0_i_67_n_0 ),
        .I1(\slvi[hmbsel][2]_INST_0_i_68_n_0 ),
        .O(hsel262_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][2]_INST_0_i_34 
       (.CI(slvi),
        .CO({hsel321_out,\slvi[hmbsel][2]_INST_0_i_34_n_1 ,\slvi[hmbsel][2]_INST_0_i_34_n_2 ,\slvi[hmbsel][2]_INST_0_i_34_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][2]_INST_0_i_69_n_0 ,\slvi[hmbsel][2]_INST_0_i_70_n_0 ,\slvi[hmbsel][2]_INST_0_i_71_n_0 ,\slvi[hmbsel][2]_INST_0_i_72_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_35 
       (.I0(\slvo[7][hconfig][6] [14]),
        .I1(\slvo[7][hconfig][6] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[7][hconfig][6] [15]),
        .I4(\slvo[7][hconfig][6] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hmbsel][2]_INST_0_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_36 
       (.I0(\slvo[7][hconfig][6] [11]),
        .I1(\slvo[7][hconfig][6] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[7][hconfig][6] [12]),
        .I4(\slvo[7][hconfig][6] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hmbsel][2]_INST_0_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_37 
       (.I0(\slvo[7][hconfig][6] [8]),
        .I1(\slvo[7][hconfig][6] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[7][hconfig][6] [9]),
        .I4(\slvo[7][hconfig][6] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hmbsel][2]_INST_0_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_38 
       (.I0(\slvo[7][hconfig][6] [5]),
        .I1(\slvo[7][hconfig][6] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[7][hconfig][6] [6]),
        .I4(\slvo[7][hconfig][6] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hmbsel][2]_INST_0_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_39 
       (.I0(\slvo[7][hconfig][6] [14]),
        .I1(\slvo[7][hconfig][6] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[7][hconfig][6] [15]),
        .I4(\slvo[7][hconfig][6] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hmbsel][2]_INST_0_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \slvi[hmbsel][2]_INST_0_i_4 
       (.I0(\slvi[hsel][2]_INST_0_i_4_n_0 ),
        .I1(\slvo[0][hconfig][6] [1]),
        .I2(\slvi[hmbsel][2]_INST_0_i_13_n_0 ),
        .I3(\slvi[hmbsel][2]_INST_0_i_14_n_0 ),
        .I4(\slvo[1][hconfig][6] [1]),
        .I5(\slvi[hsel][3]_INST_0_i_2_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_40 
       (.I0(\slvo[7][hconfig][6] [11]),
        .I1(\slvo[7][hconfig][6] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[7][hconfig][6] [12]),
        .I4(\slvo[7][hconfig][6] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hmbsel][2]_INST_0_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_41 
       (.I0(\slvo[7][hconfig][6] [8]),
        .I1(\slvo[7][hconfig][6] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[7][hconfig][6] [9]),
        .I4(\slvo[7][hconfig][6] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hmbsel][2]_INST_0_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_42 
       (.I0(\slvo[7][hconfig][6] [5]),
        .I1(\slvo[7][hconfig][6] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[7][hconfig][6] [6]),
        .I4(\slvo[7][hconfig][6] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hmbsel][2]_INST_0_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_43 
       (.I0(\slvo[6][hconfig][6] [13]),
        .I1(\slvo[6][hconfig][6] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hmbsel][2]_INST_0_i_73_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_44 
       (.I0(\slvo[6][hconfig][6] [10]),
        .I1(\slvo[6][hconfig][6] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hmbsel][2]_INST_0_i_74_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_45 
       (.I0(\slvo[6][hconfig][6] [7]),
        .I1(\slvo[6][hconfig][6] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hmbsel][2]_INST_0_i_75_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_46 
       (.I0(\slvo[6][hconfig][6] [4]),
        .I1(\slvo[6][hconfig][6] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hmbsel][2]_INST_0_i_76_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][2]_INST_0_i_47 
       (.I0(\slvo[6][hconfig][6] [9]),
        .I1(\slvo[6][hconfig][6] [7]),
        .I2(\slvo[6][hconfig][6] [8]),
        .I3(\slvo[6][hconfig][6] [4]),
        .I4(\slvo[6][hconfig][6] [5]),
        .I5(\slvo[6][hconfig][6] [6]),
        .O(\slvi[hmbsel][2]_INST_0_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][2]_INST_0_i_48 
       (.I0(\slvo[6][hconfig][6] [14]),
        .I1(\slvo[6][hconfig][6] [13]),
        .I2(\slvo[6][hconfig][6] [15]),
        .I3(\slvo[6][hconfig][6] [10]),
        .I4(\slvo[6][hconfig][6] [11]),
        .I5(\slvo[6][hconfig][6] [12]),
        .O(\slvi[hmbsel][2]_INST_0_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_49 
       (.I0(\slvo[6][hconfig][6] [13]),
        .I1(\slvo[6][hconfig][6] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hmbsel][2]_INST_0_i_77_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \slvi[hmbsel][2]_INST_0_i_5 
       (.I0(\slvi[hmbsel][2]_INST_0_i_15_n_0 ),
        .I1(\slvo[5][hconfig][6] [1]),
        .O(\slvi[hmbsel][2]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_50 
       (.I0(\slvo[6][hconfig][6] [10]),
        .I1(\slvo[6][hconfig][6] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hmbsel][2]_INST_0_i_78_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_51 
       (.I0(\slvo[6][hconfig][6] [7]),
        .I1(\slvo[6][hconfig][6] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hmbsel][2]_INST_0_i_79_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_51_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_52 
       (.I0(\slvo[6][hconfig][6] [4]),
        .I1(\slvo[6][hconfig][6] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hmbsel][2]_INST_0_i_80_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_52_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_53 
       (.I0(\slvo[4][hconfig][6] [13]),
        .I1(\slvo[4][hconfig][6] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hmbsel][2]_INST_0_i_81_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_53_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_54 
       (.I0(\slvo[4][hconfig][6] [10]),
        .I1(\slvo[4][hconfig][6] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hmbsel][2]_INST_0_i_82_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_54_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_55 
       (.I0(\slvo[4][hconfig][6] [7]),
        .I1(\slvo[4][hconfig][6] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hmbsel][2]_INST_0_i_83_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_55_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_56 
       (.I0(\slvo[4][hconfig][6] [4]),
        .I1(\slvo[4][hconfig][6] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hmbsel][2]_INST_0_i_84_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_56_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][2]_INST_0_i_57 
       (.I0(\slvo[4][hconfig][6] [9]),
        .I1(\slvo[4][hconfig][6] [7]),
        .I2(\slvo[4][hconfig][6] [8]),
        .I3(\slvo[4][hconfig][6] [4]),
        .I4(\slvo[4][hconfig][6] [5]),
        .I5(\slvo[4][hconfig][6] [6]),
        .O(\slvi[hmbsel][2]_INST_0_i_57_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][2]_INST_0_i_58 
       (.I0(\slvo[4][hconfig][6] [14]),
        .I1(\slvo[4][hconfig][6] [13]),
        .I2(\slvo[4][hconfig][6] [15]),
        .I3(\slvo[4][hconfig][6] [10]),
        .I4(\slvo[4][hconfig][6] [11]),
        .I5(\slvo[4][hconfig][6] [12]),
        .O(\slvi[hmbsel][2]_INST_0_i_58_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_59 
       (.I0(\slvo[4][hconfig][6] [13]),
        .I1(\slvo[4][hconfig][6] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hmbsel][2]_INST_0_i_85_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_59_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][2]_INST_0_i_6 
       (.CI(slvi),
        .CO({hsel30_out,\slvi[hmbsel][2]_INST_0_i_6_n_1 ,\slvi[hmbsel][2]_INST_0_i_6_n_2 ,\slvi[hmbsel][2]_INST_0_i_6_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][2]_INST_0_i_16_n_0 ,\slvi[hmbsel][2]_INST_0_i_17_n_0 ,\slvi[hmbsel][2]_INST_0_i_18_n_0 ,\slvi[hmbsel][2]_INST_0_i_19_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_60 
       (.I0(\slvo[4][hconfig][6] [10]),
        .I1(\slvo[4][hconfig][6] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hmbsel][2]_INST_0_i_86_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_60_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_61 
       (.I0(\slvo[4][hconfig][6] [7]),
        .I1(\slvo[4][hconfig][6] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hmbsel][2]_INST_0_i_87_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_61_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_62 
       (.I0(\slvo[4][hconfig][6] [4]),
        .I1(\slvo[4][hconfig][6] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hmbsel][2]_INST_0_i_88_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_62_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_63 
       (.I0(\slvo[5][hconfig][6] [13]),
        .I1(\slvo[5][hconfig][6] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hmbsel][2]_INST_0_i_89_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_63_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_64 
       (.I0(\slvo[5][hconfig][6] [10]),
        .I1(\slvo[5][hconfig][6] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hmbsel][2]_INST_0_i_90_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_64_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_65 
       (.I0(\slvo[5][hconfig][6] [7]),
        .I1(\slvo[5][hconfig][6] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hmbsel][2]_INST_0_i_91_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_65_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_66 
       (.I0(\slvo[5][hconfig][6] [4]),
        .I1(\slvo[5][hconfig][6] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hmbsel][2]_INST_0_i_92_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_66_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][2]_INST_0_i_67 
       (.I0(\slvo[5][hconfig][6] [9]),
        .I1(\slvo[5][hconfig][6] [7]),
        .I2(\slvo[5][hconfig][6] [8]),
        .I3(\slvo[5][hconfig][6] [4]),
        .I4(\slvo[5][hconfig][6] [5]),
        .I5(\slvo[5][hconfig][6] [6]),
        .O(\slvi[hmbsel][2]_INST_0_i_67_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][2]_INST_0_i_68 
       (.I0(\slvo[5][hconfig][6] [14]),
        .I1(\slvo[5][hconfig][6] [13]),
        .I2(\slvo[5][hconfig][6] [15]),
        .I3(\slvo[5][hconfig][6] [10]),
        .I4(\slvo[5][hconfig][6] [11]),
        .I5(\slvo[5][hconfig][6] [12]),
        .O(\slvi[hmbsel][2]_INST_0_i_68_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_69 
       (.I0(\slvo[5][hconfig][6] [13]),
        .I1(\slvo[5][hconfig][6] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hmbsel][2]_INST_0_i_93_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_69_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][2]_INST_0_i_7 
       (.I0(\slvi[hmbsel][2]_INST_0_i_20_n_0 ),
        .I1(\slvi[hmbsel][2]_INST_0_i_21_n_0 ),
        .O(hsel221_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_70 
       (.I0(\slvo[5][hconfig][6] [10]),
        .I1(\slvo[5][hconfig][6] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hmbsel][2]_INST_0_i_94_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_70_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_71 
       (.I0(\slvo[5][hconfig][6] [7]),
        .I1(\slvo[5][hconfig][6] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hmbsel][2]_INST_0_i_95_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_71_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][2]_INST_0_i_72 
       (.I0(\slvo[5][hconfig][6] [4]),
        .I1(\slvo[5][hconfig][6] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hmbsel][2]_INST_0_i_96_n_0 ),
        .O(\slvi[hmbsel][2]_INST_0_i_72_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_73 
       (.I0(\slvo[6][hconfig][6] [14]),
        .I1(\slvo[6][hconfig][6] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[6][hconfig][6] [15]),
        .I4(\slvo[6][hconfig][6] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hmbsel][2]_INST_0_i_73_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_74 
       (.I0(\slvo[6][hconfig][6] [11]),
        .I1(\slvo[6][hconfig][6] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[6][hconfig][6] [12]),
        .I4(\slvo[6][hconfig][6] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hmbsel][2]_INST_0_i_74_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_75 
       (.I0(\slvo[6][hconfig][6] [8]),
        .I1(\slvo[6][hconfig][6] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[6][hconfig][6] [9]),
        .I4(\slvo[6][hconfig][6] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hmbsel][2]_INST_0_i_75_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_76 
       (.I0(\slvo[6][hconfig][6] [5]),
        .I1(\slvo[6][hconfig][6] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[6][hconfig][6] [6]),
        .I4(\slvo[6][hconfig][6] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hmbsel][2]_INST_0_i_76_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_77 
       (.I0(\slvo[6][hconfig][6] [14]),
        .I1(\slvo[6][hconfig][6] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[6][hconfig][6] [15]),
        .I4(\slvo[6][hconfig][6] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hmbsel][2]_INST_0_i_77_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_78 
       (.I0(\slvo[6][hconfig][6] [11]),
        .I1(\slvo[6][hconfig][6] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[6][hconfig][6] [12]),
        .I4(\slvo[6][hconfig][6] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hmbsel][2]_INST_0_i_78_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_79 
       (.I0(\slvo[6][hconfig][6] [8]),
        .I1(\slvo[6][hconfig][6] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[6][hconfig][6] [9]),
        .I4(\slvo[6][hconfig][6] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hmbsel][2]_INST_0_i_79_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][2]_INST_0_i_8 
       (.CI(slvi),
        .CO({hsel35_out,\slvi[hmbsel][2]_INST_0_i_8_n_1 ,\slvi[hmbsel][2]_INST_0_i_8_n_2 ,\slvi[hmbsel][2]_INST_0_i_8_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][2]_INST_0_i_22_n_0 ,\slvi[hmbsel][2]_INST_0_i_23_n_0 ,\slvi[hmbsel][2]_INST_0_i_24_n_0 ,\slvi[hmbsel][2]_INST_0_i_25_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_80 
       (.I0(\slvo[6][hconfig][6] [5]),
        .I1(\slvo[6][hconfig][6] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[6][hconfig][6] [6]),
        .I4(\slvo[6][hconfig][6] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hmbsel][2]_INST_0_i_80_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_81 
       (.I0(\slvo[4][hconfig][6] [14]),
        .I1(\slvo[4][hconfig][6] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[4][hconfig][6] [15]),
        .I4(\slvo[4][hconfig][6] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hmbsel][2]_INST_0_i_81_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_82 
       (.I0(\slvo[4][hconfig][6] [11]),
        .I1(\slvo[4][hconfig][6] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[4][hconfig][6] [12]),
        .I4(\slvo[4][hconfig][6] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hmbsel][2]_INST_0_i_82_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_83 
       (.I0(\slvo[4][hconfig][6] [8]),
        .I1(\slvo[4][hconfig][6] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[4][hconfig][6] [9]),
        .I4(\slvo[4][hconfig][6] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hmbsel][2]_INST_0_i_83_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_84 
       (.I0(\slvo[4][hconfig][6] [5]),
        .I1(\slvo[4][hconfig][6] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[4][hconfig][6] [6]),
        .I4(\slvo[4][hconfig][6] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hmbsel][2]_INST_0_i_84_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_85 
       (.I0(\slvo[4][hconfig][6] [14]),
        .I1(\slvo[4][hconfig][6] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[4][hconfig][6] [15]),
        .I4(\slvo[4][hconfig][6] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hmbsel][2]_INST_0_i_85_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_86 
       (.I0(\slvo[4][hconfig][6] [11]),
        .I1(\slvo[4][hconfig][6] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[4][hconfig][6] [12]),
        .I4(\slvo[4][hconfig][6] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hmbsel][2]_INST_0_i_86_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_87 
       (.I0(\slvo[4][hconfig][6] [8]),
        .I1(\slvo[4][hconfig][6] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[4][hconfig][6] [9]),
        .I4(\slvo[4][hconfig][6] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hmbsel][2]_INST_0_i_87_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_88 
       (.I0(\slvo[4][hconfig][6] [5]),
        .I1(\slvo[4][hconfig][6] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[4][hconfig][6] [6]),
        .I4(\slvo[4][hconfig][6] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hmbsel][2]_INST_0_i_88_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_89 
       (.I0(\slvo[5][hconfig][6] [14]),
        .I1(\slvo[5][hconfig][6] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[5][hconfig][6] [15]),
        .I4(\slvo[5][hconfig][6] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hmbsel][2]_INST_0_i_89_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    \slvi[hmbsel][2]_INST_0_i_9 
       (.I0(\slvi[haddr] [20]),
        .I1(\slvi[haddr] [21]),
        .I2(\slvi[haddr] [22]),
        .I3(\slvi[haddr] [23]),
        .I4(\slvi[haddr] [24]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hmbsel][2]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_90 
       (.I0(\slvo[5][hconfig][6] [11]),
        .I1(\slvo[5][hconfig][6] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[5][hconfig][6] [12]),
        .I4(\slvo[5][hconfig][6] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hmbsel][2]_INST_0_i_90_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_91 
       (.I0(\slvo[5][hconfig][6] [8]),
        .I1(\slvo[5][hconfig][6] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[5][hconfig][6] [9]),
        .I4(\slvo[5][hconfig][6] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hmbsel][2]_INST_0_i_91_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_92 
       (.I0(\slvo[5][hconfig][6] [5]),
        .I1(\slvo[5][hconfig][6] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[5][hconfig][6] [6]),
        .I4(\slvo[5][hconfig][6] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hmbsel][2]_INST_0_i_92_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_93 
       (.I0(\slvo[5][hconfig][6] [14]),
        .I1(\slvo[5][hconfig][6] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[5][hconfig][6] [15]),
        .I4(\slvo[5][hconfig][6] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hmbsel][2]_INST_0_i_93_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_94 
       (.I0(\slvo[5][hconfig][6] [11]),
        .I1(\slvo[5][hconfig][6] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[5][hconfig][6] [12]),
        .I4(\slvo[5][hconfig][6] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hmbsel][2]_INST_0_i_94_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_95 
       (.I0(\slvo[5][hconfig][6] [8]),
        .I1(\slvo[5][hconfig][6] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[5][hconfig][6] [9]),
        .I4(\slvo[5][hconfig][6] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hmbsel][2]_INST_0_i_95_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][2]_INST_0_i_96 
       (.I0(\slvo[5][hconfig][6] [5]),
        .I1(\slvo[5][hconfig][6] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[5][hconfig][6] [6]),
        .I4(\slvo[5][hconfig][6] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hmbsel][2]_INST_0_i_96_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \slvi[hmbsel][3]_INST_0 
       (.I0(\slvi[hmbsel][3]_INST_0_i_1_n_0 ),
        .I1(\slvo[6][hconfig][7] [1]),
        .I2(\slvi[hmbsel][3]_INST_0_i_2_n_0 ),
        .I3(\slvi[hmbsel][3]_INST_0_i_3_n_0 ),
        .I4(\slvo[5][hconfig][7] [1]),
        .O(\slvi[hmbsel] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFF8F8F8FFFFFFFF)) 
    \slvi[hmbsel][3]_INST_0_i_1 
       (.I0(\slvo[4][hconfig][7] [1]),
        .I1(\slvi[hmbsel][3]_INST_0_i_4_n_0 ),
        .I2(\slvi[hmbsel][3]_INST_0_i_5_n_0 ),
        .I3(\slvi[hmbsel][3]_INST_0_i_6_n_0 ),
        .I4(\slvo[3][hconfig][7] [1]),
        .I5(\slvi[hsel][7]_INST_0_i_2_n_0 ),
        .O(\slvi[hmbsel][3]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][3]_INST_0_i_10 
       (.CI(slvi),
        .CO({hsel315_out,\slvi[hmbsel][3]_INST_0_i_10_n_1 ,\slvi[hmbsel][3]_INST_0_i_10_n_2 ,\slvi[hmbsel][3]_INST_0_i_10_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][3]_INST_0_i_26_n_0 ,\slvi[hmbsel][3]_INST_0_i_27_n_0 ,\slvi[hmbsel][3]_INST_0_i_28_n_0 ,\slvi[hmbsel][3]_INST_0_i_29_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][3]_INST_0_i_11 
       (.I0(\slvi[hmbsel][3]_INST_0_i_30_n_0 ),
        .I1(\slvi[hmbsel][3]_INST_0_i_31_n_0 ),
        .O(hsel259_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][3]_INST_0_i_12 
       (.CI(slvi),
        .CO({hsel322_out,\slvi[hmbsel][3]_INST_0_i_12_n_1 ,\slvi[hmbsel][3]_INST_0_i_12_n_2 ,\slvi[hmbsel][3]_INST_0_i_12_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][3]_INST_0_i_32_n_0 ,\slvi[hmbsel][3]_INST_0_i_33_n_0 ,\slvi[hmbsel][3]_INST_0_i_34_n_0 ,\slvi[hmbsel][3]_INST_0_i_35_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8F00800080008000)) 
    \slvi[hmbsel][3]_INST_0_i_13 
       (.I0(hsel347_out),
        .I1(hsel219_in),
        .I2(\slvo[1][hconfig][7] [0]),
        .I3(hsel2139_in),
        .I4(hsel354_out),
        .I5(hsel330_in),
        .O(\slvi[hmbsel][3]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8F00800080008000)) 
    \slvi[hmbsel][3]_INST_0_i_14 
       (.I0(hsel355_out),
        .I1(hsel219_in),
        .I2(\slvo[0][hconfig][7] [0]),
        .I3(hsel2159_in),
        .I4(hsel362_out),
        .I5(hsel330_in),
        .O(\slvi[hmbsel][3]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8F00800080008000)) 
    \slvi[hmbsel][3]_INST_0_i_15 
       (.I0(hsel339_out),
        .I1(hsel219_in),
        .I2(\slvo[2][hconfig][7] [0]),
        .I3(hsel2119_in),
        .I4(hsel346_out),
        .I5(hsel330_in),
        .O(\slvi[hmbsel][3]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][3]_INST_0_i_16 
       (.I0(\slvo[6][hconfig][7] [13]),
        .I1(\slvo[6][hconfig][7] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hmbsel][3]_INST_0_i_36_n_0 ),
        .O(\slvi[hmbsel][3]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][3]_INST_0_i_17 
       (.I0(\slvo[6][hconfig][7] [10]),
        .I1(\slvo[6][hconfig][7] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hmbsel][3]_INST_0_i_37_n_0 ),
        .O(\slvi[hmbsel][3]_INST_0_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][3]_INST_0_i_18 
       (.I0(\slvo[6][hconfig][7] [7]),
        .I1(\slvo[6][hconfig][7] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hmbsel][3]_INST_0_i_38_n_0 ),
        .O(\slvi[hmbsel][3]_INST_0_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][3]_INST_0_i_19 
       (.I0(\slvo[6][hconfig][7] [4]),
        .I1(\slvo[6][hconfig][7] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hmbsel][3]_INST_0_i_39_n_0 ),
        .O(\slvi[hmbsel][3]_INST_0_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8F00800080008000)) 
    \slvi[hmbsel][3]_INST_0_i_2 
       (.I0(hsel37_out),
        .I1(hsel219_in),
        .I2(\slvo[6][hconfig][7] [0]),
        .I3(hsel239_in),
        .I4(hsel314_out),
        .I5(hsel330_in),
        .O(\slvi[hmbsel][3]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][3]_INST_0_i_20 
       (.I0(\slvo[6][hconfig][7] [9]),
        .I1(\slvo[6][hconfig][7] [7]),
        .I2(\slvo[6][hconfig][7] [8]),
        .I3(\slvo[6][hconfig][7] [4]),
        .I4(\slvo[6][hconfig][7] [5]),
        .I5(\slvo[6][hconfig][7] [6]),
        .O(\slvi[hmbsel][3]_INST_0_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][3]_INST_0_i_21 
       (.I0(\slvo[6][hconfig][7] [14]),
        .I1(\slvo[6][hconfig][7] [13]),
        .I2(\slvo[6][hconfig][7] [15]),
        .I3(\slvo[6][hconfig][7] [10]),
        .I4(\slvo[6][hconfig][7] [11]),
        .I5(\slvo[6][hconfig][7] [12]),
        .O(\slvi[hmbsel][3]_INST_0_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][3]_INST_0_i_22 
       (.I0(\slvo[6][hconfig][7] [13]),
        .I1(\slvo[6][hconfig][7] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hmbsel][3]_INST_0_i_40_n_0 ),
        .O(\slvi[hmbsel][3]_INST_0_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][3]_INST_0_i_23 
       (.I0(\slvo[6][hconfig][7] [10]),
        .I1(\slvo[6][hconfig][7] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hmbsel][3]_INST_0_i_41_n_0 ),
        .O(\slvi[hmbsel][3]_INST_0_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][3]_INST_0_i_24 
       (.I0(\slvo[6][hconfig][7] [7]),
        .I1(\slvo[6][hconfig][7] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hmbsel][3]_INST_0_i_42_n_0 ),
        .O(\slvi[hmbsel][3]_INST_0_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][3]_INST_0_i_25 
       (.I0(\slvo[6][hconfig][7] [4]),
        .I1(\slvo[6][hconfig][7] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hmbsel][3]_INST_0_i_43_n_0 ),
        .O(\slvi[hmbsel][3]_INST_0_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][3]_INST_0_i_26 
       (.I0(\slvo[5][hconfig][7] [13]),
        .I1(\slvo[5][hconfig][7] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hmbsel][3]_INST_0_i_44_n_0 ),
        .O(\slvi[hmbsel][3]_INST_0_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][3]_INST_0_i_27 
       (.I0(\slvo[5][hconfig][7] [10]),
        .I1(\slvo[5][hconfig][7] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hmbsel][3]_INST_0_i_45_n_0 ),
        .O(\slvi[hmbsel][3]_INST_0_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][3]_INST_0_i_28 
       (.I0(\slvo[5][hconfig][7] [7]),
        .I1(\slvo[5][hconfig][7] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hmbsel][3]_INST_0_i_46_n_0 ),
        .O(\slvi[hmbsel][3]_INST_0_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][3]_INST_0_i_29 
       (.I0(\slvo[5][hconfig][7] [4]),
        .I1(\slvo[5][hconfig][7] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hmbsel][3]_INST_0_i_47_n_0 ),
        .O(\slvi[hmbsel][3]_INST_0_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8F00800080008000)) 
    \slvi[hmbsel][3]_INST_0_i_3 
       (.I0(hsel315_out),
        .I1(hsel219_in),
        .I2(\slvo[5][hconfig][7] [0]),
        .I3(hsel259_in),
        .I4(hsel322_out),
        .I5(hsel330_in),
        .O(\slvi[hmbsel][3]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][3]_INST_0_i_30 
       (.I0(\slvo[5][hconfig][7] [9]),
        .I1(\slvo[5][hconfig][7] [7]),
        .I2(\slvo[5][hconfig][7] [8]),
        .I3(\slvo[5][hconfig][7] [4]),
        .I4(\slvo[5][hconfig][7] [5]),
        .I5(\slvo[5][hconfig][7] [6]),
        .O(\slvi[hmbsel][3]_INST_0_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hmbsel][3]_INST_0_i_31 
       (.I0(\slvo[5][hconfig][7] [14]),
        .I1(\slvo[5][hconfig][7] [13]),
        .I2(\slvo[5][hconfig][7] [15]),
        .I3(\slvo[5][hconfig][7] [10]),
        .I4(\slvo[5][hconfig][7] [11]),
        .I5(\slvo[5][hconfig][7] [12]),
        .O(\slvi[hmbsel][3]_INST_0_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][3]_INST_0_i_32 
       (.I0(\slvo[5][hconfig][7] [13]),
        .I1(\slvo[5][hconfig][7] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hmbsel][3]_INST_0_i_48_n_0 ),
        .O(\slvi[hmbsel][3]_INST_0_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][3]_INST_0_i_33 
       (.I0(\slvo[5][hconfig][7] [10]),
        .I1(\slvo[5][hconfig][7] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hmbsel][3]_INST_0_i_49_n_0 ),
        .O(\slvi[hmbsel][3]_INST_0_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][3]_INST_0_i_34 
       (.I0(\slvo[5][hconfig][7] [7]),
        .I1(\slvo[5][hconfig][7] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hmbsel][3]_INST_0_i_50_n_0 ),
        .O(\slvi[hmbsel][3]_INST_0_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hmbsel][3]_INST_0_i_35 
       (.I0(\slvo[5][hconfig][7] [4]),
        .I1(\slvo[5][hconfig][7] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hmbsel][3]_INST_0_i_51_n_0 ),
        .O(\slvi[hmbsel][3]_INST_0_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][3]_INST_0_i_36 
       (.I0(\slvo[6][hconfig][7] [14]),
        .I1(\slvo[6][hconfig][7] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[6][hconfig][7] [15]),
        .I4(\slvo[6][hconfig][7] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hmbsel][3]_INST_0_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][3]_INST_0_i_37 
       (.I0(\slvo[6][hconfig][7] [11]),
        .I1(\slvo[6][hconfig][7] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[6][hconfig][7] [12]),
        .I4(\slvo[6][hconfig][7] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hmbsel][3]_INST_0_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][3]_INST_0_i_38 
       (.I0(\slvo[6][hconfig][7] [8]),
        .I1(\slvo[6][hconfig][7] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[6][hconfig][7] [9]),
        .I4(\slvo[6][hconfig][7] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hmbsel][3]_INST_0_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][3]_INST_0_i_39 
       (.I0(\slvo[6][hconfig][7] [5]),
        .I1(\slvo[6][hconfig][7] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[6][hconfig][7] [6]),
        .I4(\slvo[6][hconfig][7] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hmbsel][3]_INST_0_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8F00800080008000)) 
    \slvi[hmbsel][3]_INST_0_i_4 
       (.I0(hsel323_out),
        .I1(hsel219_in),
        .I2(\slvo[4][hconfig][7] [0]),
        .I3(hsel279_in),
        .I4(hsel330_out),
        .I5(hsel330_in),
        .O(\slvi[hmbsel][3]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][3]_INST_0_i_40 
       (.I0(\slvo[6][hconfig][7] [14]),
        .I1(\slvo[6][hconfig][7] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[6][hconfig][7] [15]),
        .I4(\slvo[6][hconfig][7] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hmbsel][3]_INST_0_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][3]_INST_0_i_41 
       (.I0(\slvo[6][hconfig][7] [11]),
        .I1(\slvo[6][hconfig][7] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[6][hconfig][7] [12]),
        .I4(\slvo[6][hconfig][7] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hmbsel][3]_INST_0_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][3]_INST_0_i_42 
       (.I0(\slvo[6][hconfig][7] [8]),
        .I1(\slvo[6][hconfig][7] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[6][hconfig][7] [9]),
        .I4(\slvo[6][hconfig][7] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hmbsel][3]_INST_0_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][3]_INST_0_i_43 
       (.I0(\slvo[6][hconfig][7] [5]),
        .I1(\slvo[6][hconfig][7] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[6][hconfig][7] [6]),
        .I4(\slvo[6][hconfig][7] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hmbsel][3]_INST_0_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][3]_INST_0_i_44 
       (.I0(\slvo[5][hconfig][7] [14]),
        .I1(\slvo[5][hconfig][7] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[5][hconfig][7] [15]),
        .I4(\slvo[5][hconfig][7] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hmbsel][3]_INST_0_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][3]_INST_0_i_45 
       (.I0(\slvo[5][hconfig][7] [11]),
        .I1(\slvo[5][hconfig][7] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[5][hconfig][7] [12]),
        .I4(\slvo[5][hconfig][7] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hmbsel][3]_INST_0_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][3]_INST_0_i_46 
       (.I0(\slvo[5][hconfig][7] [8]),
        .I1(\slvo[5][hconfig][7] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[5][hconfig][7] [9]),
        .I4(\slvo[5][hconfig][7] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hmbsel][3]_INST_0_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][3]_INST_0_i_47 
       (.I0(\slvo[5][hconfig][7] [5]),
        .I1(\slvo[5][hconfig][7] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[5][hconfig][7] [6]),
        .I4(\slvo[5][hconfig][7] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hmbsel][3]_INST_0_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][3]_INST_0_i_48 
       (.I0(\slvo[5][hconfig][7] [14]),
        .I1(\slvo[5][hconfig][7] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[5][hconfig][7] [15]),
        .I4(\slvo[5][hconfig][7] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hmbsel][3]_INST_0_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][3]_INST_0_i_49 
       (.I0(\slvo[5][hconfig][7] [11]),
        .I1(\slvo[5][hconfig][7] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[5][hconfig][7] [12]),
        .I4(\slvo[5][hconfig][7] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hmbsel][3]_INST_0_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \slvi[hmbsel][3]_INST_0_i_5 
       (.I0(\slvo[1][hconfig][7] [1]),
        .I1(\slvi[hmbsel][3]_INST_0_i_13_n_0 ),
        .I2(\slvi[hmbsel][3]_INST_0_i_14_n_0 ),
        .I3(\slvo[0][hconfig][7] [1]),
        .I4(\slvi[hmbsel][3]_INST_0_i_15_n_0 ),
        .I5(\slvo[2][hconfig][7] [1]),
        .O(\slvi[hmbsel][3]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][3]_INST_0_i_50 
       (.I0(\slvo[5][hconfig][7] [8]),
        .I1(\slvo[5][hconfig][7] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[5][hconfig][7] [9]),
        .I4(\slvo[5][hconfig][7] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hmbsel][3]_INST_0_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hmbsel][3]_INST_0_i_51 
       (.I0(\slvo[5][hconfig][7] [5]),
        .I1(\slvo[5][hconfig][7] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[5][hconfig][7] [6]),
        .I4(\slvo[5][hconfig][7] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hmbsel][3]_INST_0_i_51_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8F00800080008000)) 
    \slvi[hmbsel][3]_INST_0_i_6 
       (.I0(hsel331_out),
        .I1(hsel219_in),
        .I2(\slvo[3][hconfig][7] [0]),
        .I3(hsel299_in),
        .I4(hsel338_out),
        .I5(hsel330_in),
        .O(\slvi[hmbsel][3]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][3]_INST_0_i_7 
       (.CI(slvi),
        .CO({hsel37_out,\slvi[hmbsel][3]_INST_0_i_7_n_1 ,\slvi[hmbsel][3]_INST_0_i_7_n_2 ,\slvi[hmbsel][3]_INST_0_i_7_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][3]_INST_0_i_16_n_0 ,\slvi[hmbsel][3]_INST_0_i_17_n_0 ,\slvi[hmbsel][3]_INST_0_i_18_n_0 ,\slvi[hmbsel][3]_INST_0_i_19_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hmbsel][3]_INST_0_i_8 
       (.I0(\slvi[hmbsel][3]_INST_0_i_20_n_0 ),
        .I1(\slvi[hmbsel][3]_INST_0_i_21_n_0 ),
        .O(hsel239_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hmbsel][3]_INST_0_i_9 
       (.CI(slvi),
        .CO({hsel314_out,\slvi[hmbsel][3]_INST_0_i_9_n_1 ,\slvi[hmbsel][3]_INST_0_i_9_n_2 ,\slvi[hmbsel][3]_INST_0_i_9_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hmbsel][3]_INST_0_i_22_n_0 ,\slvi[hmbsel][3]_INST_0_i_23_n_0 ,\slvi[hmbsel][3]_INST_0_i_24_n_0 ,\slvi[hmbsel][3]_INST_0_i_25_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hprot][0]_INST_0 
       (.I0(\slvi[hprot][0]_INST_0_i_1_n_0 ),
        .I1(\slvi[hprot][0]_INST_0_i_2_n_0 ),
        .O(\slvi[hprot] [0]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hprot][0]_INST_0_i_1 
       (.I0(\msto[3][hprot] [0]),
        .I1(\msto[2][hprot] [0]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][hprot] [0]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][hprot] [0]),
        .O(\slvi[hprot][0]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hprot][0]_INST_0_i_2 
       (.I0(\msto[7][hprot] [0]),
        .I1(\msto[6][hprot] [0]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][hprot] [0]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][hprot] [0]),
        .O(\slvi[hprot][0]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hprot][1]_INST_0 
       (.I0(\slvi[hprot][1]_INST_0_i_1_n_0 ),
        .I1(\slvi[hprot][1]_INST_0_i_2_n_0 ),
        .O(\slvi[hprot] [1]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hprot][1]_INST_0_i_1 
       (.I0(\msto[3][hprot] [1]),
        .I1(\msto[2][hprot] [1]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][hprot] [1]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][hprot] [1]),
        .O(\slvi[hprot][1]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hprot][1]_INST_0_i_2 
       (.I0(\msto[7][hprot] [1]),
        .I1(\msto[6][hprot] [1]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][hprot] [1]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][hprot] [1]),
        .O(\slvi[hprot][1]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hprot][2]_INST_0 
       (.I0(\slvi[hprot][2]_INST_0_i_1_n_0 ),
        .I1(\slvi[hprot][2]_INST_0_i_2_n_0 ),
        .O(\slvi[hprot] [2]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hprot][2]_INST_0_i_1 
       (.I0(\msto[3][hprot] [2]),
        .I1(\msto[2][hprot] [2]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][hprot] [2]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][hprot] [2]),
        .O(\slvi[hprot][2]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hprot][2]_INST_0_i_2 
       (.I0(\msto[7][hprot] [2]),
        .I1(\msto[6][hprot] [2]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][hprot] [2]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][hprot] [2]),
        .O(\slvi[hprot][2]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hprot][3]_INST_0 
       (.I0(\slvi[hprot][3]_INST_0_i_1_n_0 ),
        .I1(\slvi[hprot][3]_INST_0_i_2_n_0 ),
        .O(\slvi[hprot] [3]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hprot][3]_INST_0_i_1 
       (.I0(\msto[3][hprot] [3]),
        .I1(\msto[2][hprot] [3]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][hprot] [3]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][hprot] [3]),
        .O(\slvi[hprot][3]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hprot][3]_INST_0_i_2 
       (.I0(\msto[7][hprot] [3]),
        .I1(\msto[6][hprot] [3]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][hprot] [3]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][hprot] [3]),
        .O(\slvi[hprot][3]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBBBFBBB0)) 
    \slvi[hready]_INST_0 
       (.I0(\syncrregs.r_reg[hready_n_0_] ),
        .I1(\syncrregs.r_reg[htrans_n_0_][1] ),
        .I2(\syncrregs.r_reg[defslv]__0 ),
        .I3(\syncrregs.r_reg[cfgsel_n_0_] ),
        .I4(\slvi[hready]_INST_0_i_1_n_0 ),
        .O(\slvi[hready] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hready]_INST_0_i_1 
       (.I0(\slvi[hready]_INST_0_i_2_n_0 ),
        .I1(\slvi[hready]_INST_0_i_3_n_0 ),
        .O(\slvi[hready]_INST_0_i_1_n_0 ),
        .S(\syncrregs.r_reg[hslave]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hready]_INST_0_i_2 
       (.I0(\slvo[3][hready] ),
        .I1(\slvo[2][hready] ),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[1][hready] ),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[0][hready] ),
        .O(\slvi[hready]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hready]_INST_0_i_3 
       (.I0(slvo),
        .I1(\slvo[6][hready] ),
        .I2(\syncrregs.r_reg[hslave]__0 [1]),
        .I3(\slvo[5][hready] ),
        .I4(\syncrregs.r_reg[hslave]__0 [0]),
        .I5(\slvo[4][hready] ),
        .O(\slvi[hready]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000D5FFD5D5)) 
    \slvi[hsel][0]_INST_0 
       (.I0(\slvi[hsel][0]_INST_0_i_1_n_0 ),
        .I1(\slvi[hsel][0]_INST_0_i_2_n_0 ),
        .I2(\slvo[0][hconfig][7] [1]),
        .I3(\slvi[hsel][0]_INST_0_i_3_n_0 ),
        .I4(\slvo[0][hconfig][4] [1]),
        .I5(hsel1192_out),
        .O(\^slvi[hsel] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000053FF53FF53FF)) 
    \slvi[hsel][0]_INST_0_i_1 
       (.I0(hsel1166_out),
        .I1(hsel1173_out),
        .I2(\slvo[0][hconfig][5] [0]),
        .I3(\slvo[0][hconfig][5] [1]),
        .I4(\slvo[0][hconfig][6] [1]),
        .I5(\slvi[hsel][0]_INST_0_i_7_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hsel][0]_INST_0_i_10 
       (.I0(\slvi[hsel][0]_INST_0_i_28_n_0 ),
        .I1(\slvi[hsel][0]_INST_0_i_29_n_0 ),
        .O(hsel2159_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][0]_INST_0_i_11 
       (.CI(slvi),
        .CO({hsel362_out,\slvi[hsel][0]_INST_0_i_11_n_1 ,\slvi[hsel][0]_INST_0_i_11_n_2 ,\slvi[hsel][0]_INST_0_i_11_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][0]_INST_0_i_30_n_0 ,\slvi[hsel][0]_INST_0_i_31_n_0 ,\slvi[hsel][0]_INST_0_i_32_n_0 ,\slvi[hsel][0]_INST_0_i_33_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \slvi[hsel][0]_INST_0_i_12 
       (.I0(\slvi[hmbsel][2]_INST_0_i_9_n_0 ),
        .I1(\slvi[hmbsel][2]_INST_0_i_10_n_0 ),
        .O(hsel330_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][0]_INST_0_i_13 
       (.CI(slvi),
        .CO({hsel358_out,\slvi[hsel][0]_INST_0_i_13_n_1 ,\slvi[hsel][0]_INST_0_i_13_n_2 ,\slvi[hsel][0]_INST_0_i_13_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][0]_INST_0_i_34_n_0 ,\slvi[hsel][0]_INST_0_i_35_n_0 ,\slvi[hsel][0]_INST_0_i_36_n_0 ,\slvi[hsel][0]_INST_0_i_37_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hsel][0]_INST_0_i_14 
       (.I0(\slvi[hsel][0]_INST_0_i_38_n_0 ),
        .I1(\slvi[hsel][0]_INST_0_i_39_n_0 ),
        .O(hsel2168_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][0]_INST_0_i_15 
       (.CI(slvi),
        .CO({hsel359_out,\slvi[hsel][0]_INST_0_i_15_n_1 ,\slvi[hsel][0]_INST_0_i_15_n_2 ,\slvi[hsel][0]_INST_0_i_15_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][0]_INST_0_i_40_n_0 ,\slvi[hsel][0]_INST_0_i_41_n_0 ,\slvi[hsel][0]_INST_0_i_42_n_0 ,\slvi[hsel][0]_INST_0_i_43_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    \slvi[hsel][0]_INST_0_i_16 
       (.I0(hsel219_in),
        .I1(\slvi[haddr] [12]),
        .I2(\slvi[haddr] [13]),
        .I3(\slvi[haddr] [14]),
        .I4(\slvi[haddr] [15]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hsel][0]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][0]_INST_0_i_17 
       (.I0(\slvo[0][hconfig][5] [9]),
        .I1(\slvo[0][hconfig][5] [7]),
        .I2(\slvo[0][hconfig][5] [8]),
        .I3(\slvo[0][hconfig][5] [4]),
        .I4(\slvo[0][hconfig][5] [5]),
        .I5(\slvo[0][hconfig][5] [6]),
        .O(\slvi[hsel][0]_INST_0_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][0]_INST_0_i_18 
       (.I0(\slvo[0][hconfig][5] [14]),
        .I1(\slvo[0][hconfig][5] [13]),
        .I2(\slvo[0][hconfig][5] [15]),
        .I3(\slvo[0][hconfig][5] [10]),
        .I4(\slvo[0][hconfig][5] [11]),
        .I5(\slvo[0][hconfig][5] [12]),
        .O(\slvi[hsel][0]_INST_0_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][0]_INST_0_i_19 
       (.CI(slvi),
        .CO({hsel357_out,\slvi[hsel][0]_INST_0_i_19_n_1 ,\slvi[hsel][0]_INST_0_i_19_n_2 ,\slvi[hsel][0]_INST_0_i_19_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][0]_INST_0_i_44_n_0 ,\slvi[hsel][0]_INST_0_i_45_n_0 ,\slvi[hsel][0]_INST_0_i_46_n_0 ,\slvi[hsel][0]_INST_0_i_47_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h80808080F0000000)) 
    \slvi[hsel][0]_INST_0_i_2 
       (.I0(hsel355_out),
        .I1(hsel219_in),
        .I2(hsel2159_in),
        .I3(hsel362_out),
        .I4(hsel330_in),
        .I5(\slvo[0][hconfig][7] [0]),
        .O(\slvi[hsel][0]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][0]_INST_0_i_20 
       (.CI(slvi),
        .CO({hsel360_out,\slvi[hsel][0]_INST_0_i_20_n_1 ,\slvi[hsel][0]_INST_0_i_20_n_2 ,\slvi[hsel][0]_INST_0_i_20_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][0]_INST_0_i_48_n_0 ,\slvi[hsel][0]_INST_0_i_49_n_0 ,\slvi[hsel][0]_INST_0_i_50_n_0 ,\slvi[hsel][0]_INST_0_i_51_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][0]_INST_0_i_21 
       (.CI(slvi),
        .CO({hsel356_out,\slvi[hsel][0]_INST_0_i_21_n_1 ,\slvi[hsel][0]_INST_0_i_21_n_2 ,\slvi[hsel][0]_INST_0_i_21_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][0]_INST_0_i_52_n_0 ,\slvi[hsel][0]_INST_0_i_53_n_0 ,\slvi[hsel][0]_INST_0_i_54_n_0 ,\slvi[hsel][0]_INST_0_i_55_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hsel][0]_INST_0_i_22 
       (.I0(\slvi[hsel][0]_INST_0_i_56_n_0 ),
        .I1(\slvi[hsel][0]_INST_0_i_57_n_0 ),
        .O(hsel2162_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][0]_INST_0_i_23 
       (.CI(slvi),
        .CO({hsel361_out,\slvi[hsel][0]_INST_0_i_23_n_1 ,\slvi[hsel][0]_INST_0_i_23_n_2 ,\slvi[hsel][0]_INST_0_i_23_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][0]_INST_0_i_58_n_0 ,\slvi[hsel][0]_INST_0_i_59_n_0 ,\slvi[hsel][0]_INST_0_i_60_n_0 ,\slvi[hsel][0]_INST_0_i_61_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_24 
       (.I0(\slvo[0][hconfig][7] [13]),
        .I1(\slvo[0][hconfig][7] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hsel][0]_INST_0_i_62_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_25 
       (.I0(\slvo[0][hconfig][7] [10]),
        .I1(\slvo[0][hconfig][7] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hsel][0]_INST_0_i_63_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_26 
       (.I0(\slvo[0][hconfig][7] [7]),
        .I1(\slvo[0][hconfig][7] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hsel][0]_INST_0_i_64_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_27 
       (.I0(\slvo[0][hconfig][7] [4]),
        .I1(\slvo[0][hconfig][7] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hsel][0]_INST_0_i_65_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][0]_INST_0_i_28 
       (.I0(\slvo[0][hconfig][7] [9]),
        .I1(\slvo[0][hconfig][7] [7]),
        .I2(\slvo[0][hconfig][7] [8]),
        .I3(\slvo[0][hconfig][7] [4]),
        .I4(\slvo[0][hconfig][7] [5]),
        .I5(\slvo[0][hconfig][7] [6]),
        .O(\slvi[hsel][0]_INST_0_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][0]_INST_0_i_29 
       (.I0(\slvo[0][hconfig][7] [14]),
        .I1(\slvo[0][hconfig][7] [13]),
        .I2(\slvo[0][hconfig][7] [15]),
        .I3(\slvo[0][hconfig][7] [10]),
        .I4(\slvo[0][hconfig][7] [11]),
        .I5(\slvo[0][hconfig][7] [12]),
        .O(\slvi[hsel][0]_INST_0_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h70FF7FFF7FFF7FFF)) 
    \slvi[hsel][0]_INST_0_i_3 
       (.I0(hsel358_out),
        .I1(hsel219_in),
        .I2(\slvo[0][hconfig][4] [0]),
        .I3(hsel2168_in),
        .I4(hsel359_out),
        .I5(hsel330_in),
        .O(\slvi[hsel][0]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_30 
       (.I0(\slvo[0][hconfig][7] [13]),
        .I1(\slvo[0][hconfig][7] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hsel][0]_INST_0_i_66_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_31 
       (.I0(\slvo[0][hconfig][7] [10]),
        .I1(\slvo[0][hconfig][7] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hsel][0]_INST_0_i_67_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_32 
       (.I0(\slvo[0][hconfig][7] [7]),
        .I1(\slvo[0][hconfig][7] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hsel][0]_INST_0_i_68_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_33 
       (.I0(\slvo[0][hconfig][7] [4]),
        .I1(\slvo[0][hconfig][7] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hsel][0]_INST_0_i_69_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_34 
       (.I0(\slvo[0][hconfig][4] [13]),
        .I1(\slvo[0][hconfig][4] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hsel][0]_INST_0_i_70_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_35 
       (.I0(\slvo[0][hconfig][4] [10]),
        .I1(\slvo[0][hconfig][4] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hsel][0]_INST_0_i_71_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_36 
       (.I0(\slvo[0][hconfig][4] [7]),
        .I1(\slvo[0][hconfig][4] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hsel][0]_INST_0_i_72_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_37 
       (.I0(\slvo[0][hconfig][4] [4]),
        .I1(\slvo[0][hconfig][4] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hsel][0]_INST_0_i_73_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][0]_INST_0_i_38 
       (.I0(\slvo[0][hconfig][4] [9]),
        .I1(\slvo[0][hconfig][4] [7]),
        .I2(\slvo[0][hconfig][4] [8]),
        .I3(\slvo[0][hconfig][4] [4]),
        .I4(\slvo[0][hconfig][4] [5]),
        .I5(\slvo[0][hconfig][4] [6]),
        .O(\slvi[hsel][0]_INST_0_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][0]_INST_0_i_39 
       (.I0(\slvo[0][hconfig][4] [14]),
        .I1(\slvo[0][hconfig][4] [13]),
        .I2(\slvo[0][hconfig][4] [15]),
        .I3(\slvo[0][hconfig][4] [10]),
        .I4(\slvo[0][hconfig][4] [11]),
        .I5(\slvo[0][hconfig][4] [12]),
        .O(\slvi[hsel][0]_INST_0_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0080)) 
    \slvi[hsel][0]_INST_0_i_4 
       (.I0(\slvi[haddr] [18]),
        .I1(\slvi[haddr] [19]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hsel][0]_INST_0_i_16_n_0 ),
        .O(hsel1192_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_40 
       (.I0(\slvo[0][hconfig][4] [13]),
        .I1(\slvo[0][hconfig][4] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hsel][0]_INST_0_i_74_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_41 
       (.I0(\slvo[0][hconfig][4] [10]),
        .I1(\slvo[0][hconfig][4] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hsel][0]_INST_0_i_75_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_42 
       (.I0(\slvo[0][hconfig][4] [7]),
        .I1(\slvo[0][hconfig][4] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hsel][0]_INST_0_i_76_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_43 
       (.I0(\slvo[0][hconfig][4] [4]),
        .I1(\slvo[0][hconfig][4] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hsel][0]_INST_0_i_77_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_44 
       (.I0(\slvo[0][hconfig][5] [13]),
        .I1(\slvo[0][hconfig][5] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hsel][0]_INST_0_i_78_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_45 
       (.I0(\slvo[0][hconfig][5] [10]),
        .I1(\slvo[0][hconfig][5] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hsel][0]_INST_0_i_79_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_46 
       (.I0(\slvo[0][hconfig][5] [7]),
        .I1(\slvo[0][hconfig][5] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hsel][0]_INST_0_i_80_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_47 
       (.I0(\slvo[0][hconfig][5] [4]),
        .I1(\slvo[0][hconfig][5] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hsel][0]_INST_0_i_81_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_48 
       (.I0(\slvo[0][hconfig][5] [13]),
        .I1(\slvo[0][hconfig][5] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hsel][0]_INST_0_i_82_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_49 
       (.I0(\slvo[0][hconfig][5] [10]),
        .I1(\slvo[0][hconfig][5] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hsel][0]_INST_0_i_83_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h7000)) 
    \slvi[hsel][0]_INST_0_i_5 
       (.I0(\slvi[hsel][0]_INST_0_i_17_n_0 ),
        .I1(\slvi[hsel][0]_INST_0_i_18_n_0 ),
        .I2(hsel357_out),
        .I3(hsel219_in),
        .O(hsel1166_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_50 
       (.I0(\slvo[0][hconfig][5] [7]),
        .I1(\slvo[0][hconfig][5] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hsel][0]_INST_0_i_84_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_51 
       (.I0(\slvo[0][hconfig][5] [4]),
        .I1(\slvo[0][hconfig][5] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hsel][0]_INST_0_i_85_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_51_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_52 
       (.I0(\slvo[0][hconfig][6] [13]),
        .I1(\slvo[0][hconfig][6] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hsel][0]_INST_0_i_86_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_52_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_53 
       (.I0(\slvo[0][hconfig][6] [10]),
        .I1(\slvo[0][hconfig][6] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hsel][0]_INST_0_i_87_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_53_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_54 
       (.I0(\slvo[0][hconfig][6] [7]),
        .I1(\slvo[0][hconfig][6] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hsel][0]_INST_0_i_88_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_54_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_55 
       (.I0(\slvo[0][hconfig][6] [4]),
        .I1(\slvo[0][hconfig][6] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hsel][0]_INST_0_i_89_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_55_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][0]_INST_0_i_56 
       (.I0(\slvo[0][hconfig][6] [9]),
        .I1(\slvo[0][hconfig][6] [7]),
        .I2(\slvo[0][hconfig][6] [8]),
        .I3(\slvo[0][hconfig][6] [4]),
        .I4(\slvo[0][hconfig][6] [5]),
        .I5(\slvo[0][hconfig][6] [6]),
        .O(\slvi[hsel][0]_INST_0_i_56_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][0]_INST_0_i_57 
       (.I0(\slvo[0][hconfig][6] [14]),
        .I1(\slvo[0][hconfig][6] [13]),
        .I2(\slvo[0][hconfig][6] [15]),
        .I3(\slvo[0][hconfig][6] [10]),
        .I4(\slvo[0][hconfig][6] [11]),
        .I5(\slvo[0][hconfig][6] [12]),
        .O(\slvi[hsel][0]_INST_0_i_57_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_58 
       (.I0(\slvo[0][hconfig][6] [13]),
        .I1(\slvo[0][hconfig][6] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hsel][0]_INST_0_i_90_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_58_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_59 
       (.I0(\slvo[0][hconfig][6] [10]),
        .I1(\slvo[0][hconfig][6] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hsel][0]_INST_0_i_91_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_59_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h7000)) 
    \slvi[hsel][0]_INST_0_i_6 
       (.I0(\slvi[hsel][0]_INST_0_i_17_n_0 ),
        .I1(\slvi[hsel][0]_INST_0_i_18_n_0 ),
        .I2(hsel360_out),
        .I3(hsel330_in),
        .O(hsel1173_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_60 
       (.I0(\slvo[0][hconfig][6] [7]),
        .I1(\slvo[0][hconfig][6] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hsel][0]_INST_0_i_92_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_60_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][0]_INST_0_i_61 
       (.I0(\slvo[0][hconfig][6] [4]),
        .I1(\slvo[0][hconfig][6] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hsel][0]_INST_0_i_93_n_0 ),
        .O(\slvi[hsel][0]_INST_0_i_61_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_62 
       (.I0(\slvo[0][hconfig][7] [14]),
        .I1(\slvo[0][hconfig][7] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[0][hconfig][7] [15]),
        .I4(\slvo[0][hconfig][7] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hsel][0]_INST_0_i_62_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_63 
       (.I0(\slvo[0][hconfig][7] [11]),
        .I1(\slvo[0][hconfig][7] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[0][hconfig][7] [12]),
        .I4(\slvo[0][hconfig][7] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hsel][0]_INST_0_i_63_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_64 
       (.I0(\slvo[0][hconfig][7] [8]),
        .I1(\slvo[0][hconfig][7] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[0][hconfig][7] [9]),
        .I4(\slvo[0][hconfig][7] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hsel][0]_INST_0_i_64_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_65 
       (.I0(\slvo[0][hconfig][7] [5]),
        .I1(\slvo[0][hconfig][7] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[0][hconfig][7] [6]),
        .I4(\slvo[0][hconfig][7] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hsel][0]_INST_0_i_65_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_66 
       (.I0(\slvo[0][hconfig][7] [14]),
        .I1(\slvo[0][hconfig][7] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[0][hconfig][7] [15]),
        .I4(\slvo[0][hconfig][7] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hsel][0]_INST_0_i_66_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_67 
       (.I0(\slvo[0][hconfig][7] [11]),
        .I1(\slvo[0][hconfig][7] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[0][hconfig][7] [12]),
        .I4(\slvo[0][hconfig][7] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hsel][0]_INST_0_i_67_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_68 
       (.I0(\slvo[0][hconfig][7] [8]),
        .I1(\slvo[0][hconfig][7] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[0][hconfig][7] [9]),
        .I4(\slvo[0][hconfig][7] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hsel][0]_INST_0_i_68_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_69 
       (.I0(\slvo[0][hconfig][7] [5]),
        .I1(\slvo[0][hconfig][7] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[0][hconfig][7] [6]),
        .I4(\slvo[0][hconfig][7] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hsel][0]_INST_0_i_69_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h80808080F0000000)) 
    \slvi[hsel][0]_INST_0_i_7 
       (.I0(hsel356_out),
        .I1(hsel219_in),
        .I2(hsel2162_in),
        .I3(hsel361_out),
        .I4(hsel330_in),
        .I5(\slvo[0][hconfig][6] [0]),
        .O(\slvi[hsel][0]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_70 
       (.I0(\slvo[0][hconfig][4] [14]),
        .I1(\slvo[0][hconfig][4] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[0][hconfig][4] [15]),
        .I4(\slvo[0][hconfig][4] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hsel][0]_INST_0_i_70_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_71 
       (.I0(\slvo[0][hconfig][4] [11]),
        .I1(\slvo[0][hconfig][4] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[0][hconfig][4] [12]),
        .I4(\slvo[0][hconfig][4] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hsel][0]_INST_0_i_71_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_72 
       (.I0(\slvo[0][hconfig][4] [8]),
        .I1(\slvo[0][hconfig][4] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[0][hconfig][4] [9]),
        .I4(\slvo[0][hconfig][4] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hsel][0]_INST_0_i_72_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_73 
       (.I0(\slvo[0][hconfig][4] [5]),
        .I1(\slvo[0][hconfig][4] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[0][hconfig][4] [6]),
        .I4(\slvo[0][hconfig][4] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hsel][0]_INST_0_i_73_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_74 
       (.I0(\slvo[0][hconfig][4] [14]),
        .I1(\slvo[0][hconfig][4] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[0][hconfig][4] [15]),
        .I4(\slvo[0][hconfig][4] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hsel][0]_INST_0_i_74_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_75 
       (.I0(\slvo[0][hconfig][4] [11]),
        .I1(\slvo[0][hconfig][4] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[0][hconfig][4] [12]),
        .I4(\slvo[0][hconfig][4] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hsel][0]_INST_0_i_75_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_76 
       (.I0(\slvo[0][hconfig][4] [8]),
        .I1(\slvo[0][hconfig][4] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[0][hconfig][4] [9]),
        .I4(\slvo[0][hconfig][4] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hsel][0]_INST_0_i_76_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_77 
       (.I0(\slvo[0][hconfig][4] [5]),
        .I1(\slvo[0][hconfig][4] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[0][hconfig][4] [6]),
        .I4(\slvo[0][hconfig][4] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hsel][0]_INST_0_i_77_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_78 
       (.I0(\slvo[0][hconfig][5] [14]),
        .I1(\slvo[0][hconfig][5] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[0][hconfig][5] [15]),
        .I4(\slvo[0][hconfig][5] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hsel][0]_INST_0_i_78_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_79 
       (.I0(\slvo[0][hconfig][5] [11]),
        .I1(\slvo[0][hconfig][5] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[0][hconfig][5] [12]),
        .I4(\slvo[0][hconfig][5] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hsel][0]_INST_0_i_79_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][0]_INST_0_i_8 
       (.CI(slvi),
        .CO({hsel355_out,\slvi[hsel][0]_INST_0_i_8_n_1 ,\slvi[hsel][0]_INST_0_i_8_n_2 ,\slvi[hsel][0]_INST_0_i_8_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][0]_INST_0_i_24_n_0 ,\slvi[hsel][0]_INST_0_i_25_n_0 ,\slvi[hsel][0]_INST_0_i_26_n_0 ,\slvi[hsel][0]_INST_0_i_27_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_80 
       (.I0(\slvo[0][hconfig][5] [8]),
        .I1(\slvo[0][hconfig][5] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[0][hconfig][5] [9]),
        .I4(\slvo[0][hconfig][5] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hsel][0]_INST_0_i_80_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_81 
       (.I0(\slvo[0][hconfig][5] [5]),
        .I1(\slvo[0][hconfig][5] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[0][hconfig][5] [6]),
        .I4(\slvo[0][hconfig][5] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hsel][0]_INST_0_i_81_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_82 
       (.I0(\slvo[0][hconfig][5] [14]),
        .I1(\slvo[0][hconfig][5] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[0][hconfig][5] [15]),
        .I4(\slvo[0][hconfig][5] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hsel][0]_INST_0_i_82_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_83 
       (.I0(\slvo[0][hconfig][5] [11]),
        .I1(\slvo[0][hconfig][5] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[0][hconfig][5] [12]),
        .I4(\slvo[0][hconfig][5] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hsel][0]_INST_0_i_83_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_84 
       (.I0(\slvo[0][hconfig][5] [8]),
        .I1(\slvo[0][hconfig][5] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[0][hconfig][5] [9]),
        .I4(\slvo[0][hconfig][5] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hsel][0]_INST_0_i_84_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_85 
       (.I0(\slvo[0][hconfig][5] [5]),
        .I1(\slvo[0][hconfig][5] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[0][hconfig][5] [6]),
        .I4(\slvo[0][hconfig][5] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hsel][0]_INST_0_i_85_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_86 
       (.I0(\slvo[0][hconfig][6] [14]),
        .I1(\slvo[0][hconfig][6] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[0][hconfig][6] [15]),
        .I4(\slvo[0][hconfig][6] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hsel][0]_INST_0_i_86_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_87 
       (.I0(\slvo[0][hconfig][6] [11]),
        .I1(\slvo[0][hconfig][6] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[0][hconfig][6] [12]),
        .I4(\slvo[0][hconfig][6] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hsel][0]_INST_0_i_87_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_88 
       (.I0(\slvo[0][hconfig][6] [8]),
        .I1(\slvo[0][hconfig][6] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[0][hconfig][6] [9]),
        .I4(\slvo[0][hconfig][6] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hsel][0]_INST_0_i_88_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_89 
       (.I0(\slvo[0][hconfig][6] [5]),
        .I1(\slvo[0][hconfig][6] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[0][hconfig][6] [6]),
        .I4(\slvo[0][hconfig][6] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hsel][0]_INST_0_i_89_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \slvi[hsel][0]_INST_0_i_9 
       (.I0(\slvi[hmbsel][2]_INST_0_i_10_n_0 ),
        .I1(\slvi[hmbsel][2]_INST_0_i_9_n_0 ),
        .O(hsel219_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_90 
       (.I0(\slvo[0][hconfig][6] [14]),
        .I1(\slvo[0][hconfig][6] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[0][hconfig][6] [15]),
        .I4(\slvo[0][hconfig][6] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hsel][0]_INST_0_i_90_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_91 
       (.I0(\slvo[0][hconfig][6] [11]),
        .I1(\slvo[0][hconfig][6] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[0][hconfig][6] [12]),
        .I4(\slvo[0][hconfig][6] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hsel][0]_INST_0_i_91_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_92 
       (.I0(\slvo[0][hconfig][6] [8]),
        .I1(\slvo[0][hconfig][6] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[0][hconfig][6] [9]),
        .I4(\slvo[0][hconfig][6] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hsel][0]_INST_0_i_92_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][0]_INST_0_i_93 
       (.I0(\slvo[0][hconfig][6] [5]),
        .I1(\slvo[0][hconfig][6] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[0][hconfig][6] [6]),
        .I4(\slvo[0][hconfig][6] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hsel][0]_INST_0_i_93_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \slvi[hsel][1]_INST_0 
       (.I0(\slvi[hsel][1]_INST_0_i_1_n_0 ),
        .I1(hsel1192_out),
        .O(\^slvi[hsel] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF777F777F777)) 
    \slvi[hsel][1]_INST_0_i_1 
       (.I0(\slvi[hsel][1]_INST_0_i_2_n_0 ),
        .I1(\slvi[hsel][1]_INST_0_i_3_n_0 ),
        .I2(\slvo[1][hconfig][7] [1]),
        .I3(\slvi[hsel][1]_INST_0_i_4_n_0 ),
        .I4(\slvi[hsel][1]_INST_0_i_5_n_0 ),
        .I5(\slvo[1][hconfig][6] [1]),
        .O(\slvi[hsel][1]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][1]_INST_0_i_10 
       (.CI(slvi),
        .CO({hsel354_out,\slvi[hsel][1]_INST_0_i_10_n_1 ,\slvi[hsel][1]_INST_0_i_10_n_2 ,\slvi[hsel][1]_INST_0_i_10_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][1]_INST_0_i_26_n_0 ,\slvi[hsel][1]_INST_0_i_27_n_0 ,\slvi[hsel][1]_INST_0_i_28_n_0 ,\slvi[hsel][1]_INST_0_i_29_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][1]_INST_0_i_11 
       (.CI(slvi),
        .CO({hsel348_out,\slvi[hsel][1]_INST_0_i_11_n_1 ,\slvi[hsel][1]_INST_0_i_11_n_2 ,\slvi[hsel][1]_INST_0_i_11_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][1]_INST_0_i_30_n_0 ,\slvi[hsel][1]_INST_0_i_31_n_0 ,\slvi[hsel][1]_INST_0_i_32_n_0 ,\slvi[hsel][1]_INST_0_i_33_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hsel][1]_INST_0_i_12 
       (.I0(\slvi[hsel][1]_INST_0_i_34_n_0 ),
        .I1(\slvi[hsel][1]_INST_0_i_35_n_0 ),
        .O(hsel2142_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][1]_INST_0_i_13 
       (.CI(slvi),
        .CO({hsel353_out,\slvi[hsel][1]_INST_0_i_13_n_1 ,\slvi[hsel][1]_INST_0_i_13_n_2 ,\slvi[hsel][1]_INST_0_i_13_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][1]_INST_0_i_36_n_0 ,\slvi[hsel][1]_INST_0_i_37_n_0 ,\slvi[hsel][1]_INST_0_i_38_n_0 ,\slvi[hsel][1]_INST_0_i_39_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][1]_INST_0_i_14 
       (.CI(slvi),
        .CO({hsel350_out,\slvi[hsel][1]_INST_0_i_14_n_1 ,\slvi[hsel][1]_INST_0_i_14_n_2 ,\slvi[hsel][1]_INST_0_i_14_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][1]_INST_0_i_40_n_0 ,\slvi[hsel][1]_INST_0_i_41_n_0 ,\slvi[hsel][1]_INST_0_i_42_n_0 ,\slvi[hsel][1]_INST_0_i_43_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hsel][1]_INST_0_i_15 
       (.I0(\slvi[hsel][1]_INST_0_i_44_n_0 ),
        .I1(\slvi[hsel][1]_INST_0_i_45_n_0 ),
        .O(hsel2148_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][1]_INST_0_i_16 
       (.CI(slvi),
        .CO({hsel351_out,\slvi[hsel][1]_INST_0_i_16_n_1 ,\slvi[hsel][1]_INST_0_i_16_n_2 ,\slvi[hsel][1]_INST_0_i_16_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][1]_INST_0_i_46_n_0 ,\slvi[hsel][1]_INST_0_i_47_n_0 ,\slvi[hsel][1]_INST_0_i_48_n_0 ,\slvi[hsel][1]_INST_0_i_49_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][1]_INST_0_i_17 
       (.CI(slvi),
        .CO({hsel349_out,\slvi[hsel][1]_INST_0_i_17_n_1 ,\slvi[hsel][1]_INST_0_i_17_n_2 ,\slvi[hsel][1]_INST_0_i_17_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][1]_INST_0_i_50_n_0 ,\slvi[hsel][1]_INST_0_i_51_n_0 ,\slvi[hsel][1]_INST_0_i_52_n_0 ,\slvi[hsel][1]_INST_0_i_53_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hsel][1]_INST_0_i_18 
       (.I0(\slvi[hsel][1]_INST_0_i_54_n_0 ),
        .I1(\slvi[hsel][1]_INST_0_i_55_n_0 ),
        .O(hsel2145_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][1]_INST_0_i_19 
       (.CI(slvi),
        .CO({hsel352_out,\slvi[hsel][1]_INST_0_i_19_n_1 ,\slvi[hsel][1]_INST_0_i_19_n_2 ,\slvi[hsel][1]_INST_0_i_19_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][1]_INST_0_i_56_n_0 ,\slvi[hsel][1]_INST_0_i_57_n_0 ,\slvi[hsel][1]_INST_0_i_58_n_0 ,\slvi[hsel][1]_INST_0_i_59_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hsel][1]_INST_0_i_2 
       (.I0(\slvo[1][hconfig][4] [1]),
        .I1(\slvi[hsel][1]_INST_0_i_6_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_20 
       (.I0(\slvo[1][hconfig][7] [13]),
        .I1(\slvo[1][hconfig][7] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hsel][1]_INST_0_i_60_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_21 
       (.I0(\slvo[1][hconfig][7] [10]),
        .I1(\slvo[1][hconfig][7] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hsel][1]_INST_0_i_61_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_22 
       (.I0(\slvo[1][hconfig][7] [7]),
        .I1(\slvo[1][hconfig][7] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hsel][1]_INST_0_i_62_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_23 
       (.I0(\slvo[1][hconfig][7] [4]),
        .I1(\slvo[1][hconfig][7] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hsel][1]_INST_0_i_63_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][1]_INST_0_i_24 
       (.I0(\slvo[1][hconfig][7] [9]),
        .I1(\slvo[1][hconfig][7] [7]),
        .I2(\slvo[1][hconfig][7] [8]),
        .I3(\slvo[1][hconfig][7] [4]),
        .I4(\slvo[1][hconfig][7] [5]),
        .I5(\slvo[1][hconfig][7] [6]),
        .O(\slvi[hsel][1]_INST_0_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][1]_INST_0_i_25 
       (.I0(\slvo[1][hconfig][7] [14]),
        .I1(\slvo[1][hconfig][7] [13]),
        .I2(\slvo[1][hconfig][7] [15]),
        .I3(\slvo[1][hconfig][7] [10]),
        .I4(\slvo[1][hconfig][7] [11]),
        .I5(\slvo[1][hconfig][7] [12]),
        .O(\slvi[hsel][1]_INST_0_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_26 
       (.I0(\slvo[1][hconfig][7] [13]),
        .I1(\slvo[1][hconfig][7] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hsel][1]_INST_0_i_64_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_27 
       (.I0(\slvo[1][hconfig][7] [10]),
        .I1(\slvo[1][hconfig][7] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hsel][1]_INST_0_i_65_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_28 
       (.I0(\slvo[1][hconfig][7] [7]),
        .I1(\slvo[1][hconfig][7] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hsel][1]_INST_0_i_66_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_29 
       (.I0(\slvo[1][hconfig][7] [4]),
        .I1(\slvo[1][hconfig][7] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hsel][1]_INST_0_i_67_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hsel][1]_INST_0_i_3 
       (.I0(\slvo[1][hconfig][5] [1]),
        .I1(\slvi[hsel][1]_INST_0_i_7_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_30 
       (.I0(\slvo[1][hconfig][6] [13]),
        .I1(\slvo[1][hconfig][6] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hsel][1]_INST_0_i_68_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_31 
       (.I0(\slvo[1][hconfig][6] [10]),
        .I1(\slvo[1][hconfig][6] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hsel][1]_INST_0_i_69_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_32 
       (.I0(\slvo[1][hconfig][6] [7]),
        .I1(\slvo[1][hconfig][6] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hsel][1]_INST_0_i_70_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_33 
       (.I0(\slvo[1][hconfig][6] [4]),
        .I1(\slvo[1][hconfig][6] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hsel][1]_INST_0_i_71_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][1]_INST_0_i_34 
       (.I0(\slvo[1][hconfig][6] [9]),
        .I1(\slvo[1][hconfig][6] [7]),
        .I2(\slvo[1][hconfig][6] [8]),
        .I3(\slvo[1][hconfig][6] [4]),
        .I4(\slvo[1][hconfig][6] [5]),
        .I5(\slvo[1][hconfig][6] [6]),
        .O(\slvi[hsel][1]_INST_0_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][1]_INST_0_i_35 
       (.I0(\slvo[1][hconfig][6] [14]),
        .I1(\slvo[1][hconfig][6] [13]),
        .I2(\slvo[1][hconfig][6] [15]),
        .I3(\slvo[1][hconfig][6] [10]),
        .I4(\slvo[1][hconfig][6] [11]),
        .I5(\slvo[1][hconfig][6] [12]),
        .O(\slvi[hsel][1]_INST_0_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_36 
       (.I0(\slvo[1][hconfig][6] [13]),
        .I1(\slvo[1][hconfig][6] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hsel][1]_INST_0_i_72_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_37 
       (.I0(\slvo[1][hconfig][6] [10]),
        .I1(\slvo[1][hconfig][6] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hsel][1]_INST_0_i_73_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_38 
       (.I0(\slvo[1][hconfig][6] [7]),
        .I1(\slvo[1][hconfig][6] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hsel][1]_INST_0_i_74_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_39 
       (.I0(\slvo[1][hconfig][6] [4]),
        .I1(\slvo[1][hconfig][6] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hsel][1]_INST_0_i_75_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h80808080F0000000)) 
    \slvi[hsel][1]_INST_0_i_4 
       (.I0(hsel347_out),
        .I1(hsel219_in),
        .I2(hsel2139_in),
        .I3(hsel354_out),
        .I4(hsel330_in),
        .I5(\slvo[1][hconfig][7] [0]),
        .O(\slvi[hsel][1]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_40 
       (.I0(\slvo[1][hconfig][4] [13]),
        .I1(\slvo[1][hconfig][4] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hsel][1]_INST_0_i_76_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_41 
       (.I0(\slvo[1][hconfig][4] [10]),
        .I1(\slvo[1][hconfig][4] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hsel][1]_INST_0_i_77_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_42 
       (.I0(\slvo[1][hconfig][4] [7]),
        .I1(\slvo[1][hconfig][4] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hsel][1]_INST_0_i_78_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_43 
       (.I0(\slvo[1][hconfig][4] [4]),
        .I1(\slvo[1][hconfig][4] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hsel][1]_INST_0_i_79_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][1]_INST_0_i_44 
       (.I0(\slvo[1][hconfig][4] [9]),
        .I1(\slvo[1][hconfig][4] [7]),
        .I2(\slvo[1][hconfig][4] [8]),
        .I3(\slvo[1][hconfig][4] [4]),
        .I4(\slvo[1][hconfig][4] [5]),
        .I5(\slvo[1][hconfig][4] [6]),
        .O(\slvi[hsel][1]_INST_0_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][1]_INST_0_i_45 
       (.I0(\slvo[1][hconfig][4] [14]),
        .I1(\slvo[1][hconfig][4] [13]),
        .I2(\slvo[1][hconfig][4] [15]),
        .I3(\slvo[1][hconfig][4] [10]),
        .I4(\slvo[1][hconfig][4] [11]),
        .I5(\slvo[1][hconfig][4] [12]),
        .O(\slvi[hsel][1]_INST_0_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_46 
       (.I0(\slvo[1][hconfig][4] [13]),
        .I1(\slvo[1][hconfig][4] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hsel][1]_INST_0_i_80_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_47 
       (.I0(\slvo[1][hconfig][4] [10]),
        .I1(\slvo[1][hconfig][4] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hsel][1]_INST_0_i_81_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_48 
       (.I0(\slvo[1][hconfig][4] [7]),
        .I1(\slvo[1][hconfig][4] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hsel][1]_INST_0_i_82_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_49 
       (.I0(\slvo[1][hconfig][4] [4]),
        .I1(\slvo[1][hconfig][4] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hsel][1]_INST_0_i_83_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h80808080F0000000)) 
    \slvi[hsel][1]_INST_0_i_5 
       (.I0(hsel348_out),
        .I1(hsel219_in),
        .I2(hsel2142_in),
        .I3(hsel353_out),
        .I4(hsel330_in),
        .I5(\slvo[1][hconfig][6] [0]),
        .O(\slvi[hsel][1]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_50 
       (.I0(\slvo[1][hconfig][5] [13]),
        .I1(\slvo[1][hconfig][5] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hsel][1]_INST_0_i_84_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_51 
       (.I0(\slvo[1][hconfig][5] [10]),
        .I1(\slvo[1][hconfig][5] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hsel][1]_INST_0_i_85_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_51_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_52 
       (.I0(\slvo[1][hconfig][5] [7]),
        .I1(\slvo[1][hconfig][5] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hsel][1]_INST_0_i_86_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_52_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_53 
       (.I0(\slvo[1][hconfig][5] [4]),
        .I1(\slvo[1][hconfig][5] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hsel][1]_INST_0_i_87_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_53_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][1]_INST_0_i_54 
       (.I0(\slvo[1][hconfig][5] [9]),
        .I1(\slvo[1][hconfig][5] [7]),
        .I2(\slvo[1][hconfig][5] [8]),
        .I3(\slvo[1][hconfig][5] [4]),
        .I4(\slvo[1][hconfig][5] [5]),
        .I5(\slvo[1][hconfig][5] [6]),
        .O(\slvi[hsel][1]_INST_0_i_54_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][1]_INST_0_i_55 
       (.I0(\slvo[1][hconfig][5] [14]),
        .I1(\slvo[1][hconfig][5] [13]),
        .I2(\slvo[1][hconfig][5] [15]),
        .I3(\slvo[1][hconfig][5] [10]),
        .I4(\slvo[1][hconfig][5] [11]),
        .I5(\slvo[1][hconfig][5] [12]),
        .O(\slvi[hsel][1]_INST_0_i_55_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_56 
       (.I0(\slvo[1][hconfig][5] [13]),
        .I1(\slvo[1][hconfig][5] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hsel][1]_INST_0_i_88_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_56_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_57 
       (.I0(\slvo[1][hconfig][5] [10]),
        .I1(\slvo[1][hconfig][5] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hsel][1]_INST_0_i_89_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_57_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_58 
       (.I0(\slvo[1][hconfig][5] [7]),
        .I1(\slvo[1][hconfig][5] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hsel][1]_INST_0_i_90_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_58_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][1]_INST_0_i_59 
       (.I0(\slvo[1][hconfig][5] [4]),
        .I1(\slvo[1][hconfig][5] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hsel][1]_INST_0_i_91_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_59_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000808030003000)) 
    \slvi[hsel][1]_INST_0_i_6 
       (.I0(hsel350_out),
        .I1(\slvo[1][hconfig][4] [0]),
        .I2(hsel2148_in),
        .I3(hsel351_out),
        .I4(\slvi[hmbsel][2]_INST_0_i_9_n_0 ),
        .I5(\slvi[hmbsel][2]_INST_0_i_10_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_60 
       (.I0(\slvo[1][hconfig][7] [14]),
        .I1(\slvo[1][hconfig][7] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[1][hconfig][7] [15]),
        .I4(\slvo[1][hconfig][7] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hsel][1]_INST_0_i_60_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_61 
       (.I0(\slvo[1][hconfig][7] [11]),
        .I1(\slvo[1][hconfig][7] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[1][hconfig][7] [12]),
        .I4(\slvo[1][hconfig][7] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hsel][1]_INST_0_i_61_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_62 
       (.I0(\slvo[1][hconfig][7] [8]),
        .I1(\slvo[1][hconfig][7] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[1][hconfig][7] [9]),
        .I4(\slvo[1][hconfig][7] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hsel][1]_INST_0_i_62_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_63 
       (.I0(\slvo[1][hconfig][7] [5]),
        .I1(\slvo[1][hconfig][7] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[1][hconfig][7] [6]),
        .I4(\slvo[1][hconfig][7] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hsel][1]_INST_0_i_63_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_64 
       (.I0(\slvo[1][hconfig][7] [14]),
        .I1(\slvo[1][hconfig][7] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[1][hconfig][7] [15]),
        .I4(\slvo[1][hconfig][7] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hsel][1]_INST_0_i_64_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_65 
       (.I0(\slvo[1][hconfig][7] [11]),
        .I1(\slvo[1][hconfig][7] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[1][hconfig][7] [12]),
        .I4(\slvo[1][hconfig][7] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hsel][1]_INST_0_i_65_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_66 
       (.I0(\slvo[1][hconfig][7] [8]),
        .I1(\slvo[1][hconfig][7] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[1][hconfig][7] [9]),
        .I4(\slvo[1][hconfig][7] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hsel][1]_INST_0_i_66_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_67 
       (.I0(\slvo[1][hconfig][7] [5]),
        .I1(\slvo[1][hconfig][7] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[1][hconfig][7] [6]),
        .I4(\slvo[1][hconfig][7] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hsel][1]_INST_0_i_67_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_68 
       (.I0(\slvo[1][hconfig][6] [14]),
        .I1(\slvo[1][hconfig][6] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[1][hconfig][6] [15]),
        .I4(\slvo[1][hconfig][6] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hsel][1]_INST_0_i_68_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_69 
       (.I0(\slvo[1][hconfig][6] [11]),
        .I1(\slvo[1][hconfig][6] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[1][hconfig][6] [12]),
        .I4(\slvo[1][hconfig][6] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hsel][1]_INST_0_i_69_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000808030003000)) 
    \slvi[hsel][1]_INST_0_i_7 
       (.I0(hsel349_out),
        .I1(\slvo[1][hconfig][5] [0]),
        .I2(hsel2145_in),
        .I3(hsel352_out),
        .I4(\slvi[hmbsel][2]_INST_0_i_9_n_0 ),
        .I5(\slvi[hmbsel][2]_INST_0_i_10_n_0 ),
        .O(\slvi[hsel][1]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_70 
       (.I0(\slvo[1][hconfig][6] [8]),
        .I1(\slvo[1][hconfig][6] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[1][hconfig][6] [9]),
        .I4(\slvo[1][hconfig][6] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hsel][1]_INST_0_i_70_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_71 
       (.I0(\slvo[1][hconfig][6] [5]),
        .I1(\slvo[1][hconfig][6] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[1][hconfig][6] [6]),
        .I4(\slvo[1][hconfig][6] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hsel][1]_INST_0_i_71_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_72 
       (.I0(\slvo[1][hconfig][6] [14]),
        .I1(\slvo[1][hconfig][6] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[1][hconfig][6] [15]),
        .I4(\slvo[1][hconfig][6] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hsel][1]_INST_0_i_72_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_73 
       (.I0(\slvo[1][hconfig][6] [11]),
        .I1(\slvo[1][hconfig][6] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[1][hconfig][6] [12]),
        .I4(\slvo[1][hconfig][6] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hsel][1]_INST_0_i_73_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_74 
       (.I0(\slvo[1][hconfig][6] [8]),
        .I1(\slvo[1][hconfig][6] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[1][hconfig][6] [9]),
        .I4(\slvo[1][hconfig][6] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hsel][1]_INST_0_i_74_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_75 
       (.I0(\slvo[1][hconfig][6] [5]),
        .I1(\slvo[1][hconfig][6] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[1][hconfig][6] [6]),
        .I4(\slvo[1][hconfig][6] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hsel][1]_INST_0_i_75_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_76 
       (.I0(\slvo[1][hconfig][4] [14]),
        .I1(\slvo[1][hconfig][4] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[1][hconfig][4] [15]),
        .I4(\slvo[1][hconfig][4] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hsel][1]_INST_0_i_76_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_77 
       (.I0(\slvo[1][hconfig][4] [11]),
        .I1(\slvo[1][hconfig][4] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[1][hconfig][4] [12]),
        .I4(\slvo[1][hconfig][4] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hsel][1]_INST_0_i_77_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_78 
       (.I0(\slvo[1][hconfig][4] [8]),
        .I1(\slvo[1][hconfig][4] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[1][hconfig][4] [9]),
        .I4(\slvo[1][hconfig][4] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hsel][1]_INST_0_i_78_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_79 
       (.I0(\slvo[1][hconfig][4] [5]),
        .I1(\slvo[1][hconfig][4] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[1][hconfig][4] [6]),
        .I4(\slvo[1][hconfig][4] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hsel][1]_INST_0_i_79_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][1]_INST_0_i_8 
       (.CI(slvi),
        .CO({hsel347_out,\slvi[hsel][1]_INST_0_i_8_n_1 ,\slvi[hsel][1]_INST_0_i_8_n_2 ,\slvi[hsel][1]_INST_0_i_8_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][1]_INST_0_i_20_n_0 ,\slvi[hsel][1]_INST_0_i_21_n_0 ,\slvi[hsel][1]_INST_0_i_22_n_0 ,\slvi[hsel][1]_INST_0_i_23_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_80 
       (.I0(\slvo[1][hconfig][4] [14]),
        .I1(\slvo[1][hconfig][4] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[1][hconfig][4] [15]),
        .I4(\slvo[1][hconfig][4] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hsel][1]_INST_0_i_80_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_81 
       (.I0(\slvo[1][hconfig][4] [11]),
        .I1(\slvo[1][hconfig][4] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[1][hconfig][4] [12]),
        .I4(\slvo[1][hconfig][4] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hsel][1]_INST_0_i_81_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_82 
       (.I0(\slvo[1][hconfig][4] [8]),
        .I1(\slvo[1][hconfig][4] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[1][hconfig][4] [9]),
        .I4(\slvo[1][hconfig][4] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hsel][1]_INST_0_i_82_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_83 
       (.I0(\slvo[1][hconfig][4] [5]),
        .I1(\slvo[1][hconfig][4] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[1][hconfig][4] [6]),
        .I4(\slvo[1][hconfig][4] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hsel][1]_INST_0_i_83_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_84 
       (.I0(\slvo[1][hconfig][5] [14]),
        .I1(\slvo[1][hconfig][5] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[1][hconfig][5] [15]),
        .I4(\slvo[1][hconfig][5] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hsel][1]_INST_0_i_84_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_85 
       (.I0(\slvo[1][hconfig][5] [11]),
        .I1(\slvo[1][hconfig][5] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[1][hconfig][5] [12]),
        .I4(\slvo[1][hconfig][5] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hsel][1]_INST_0_i_85_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_86 
       (.I0(\slvo[1][hconfig][5] [8]),
        .I1(\slvo[1][hconfig][5] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[1][hconfig][5] [9]),
        .I4(\slvo[1][hconfig][5] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hsel][1]_INST_0_i_86_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_87 
       (.I0(\slvo[1][hconfig][5] [5]),
        .I1(\slvo[1][hconfig][5] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[1][hconfig][5] [6]),
        .I4(\slvo[1][hconfig][5] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hsel][1]_INST_0_i_87_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_88 
       (.I0(\slvo[1][hconfig][5] [14]),
        .I1(\slvo[1][hconfig][5] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[1][hconfig][5] [15]),
        .I4(\slvo[1][hconfig][5] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hsel][1]_INST_0_i_88_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_89 
       (.I0(\slvo[1][hconfig][5] [11]),
        .I1(\slvo[1][hconfig][5] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[1][hconfig][5] [12]),
        .I4(\slvo[1][hconfig][5] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hsel][1]_INST_0_i_89_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hsel][1]_INST_0_i_9 
       (.I0(\slvi[hsel][1]_INST_0_i_24_n_0 ),
        .I1(\slvi[hsel][1]_INST_0_i_25_n_0 ),
        .O(hsel2139_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_90 
       (.I0(\slvo[1][hconfig][5] [8]),
        .I1(\slvo[1][hconfig][5] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[1][hconfig][5] [9]),
        .I4(\slvo[1][hconfig][5] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hsel][1]_INST_0_i_90_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][1]_INST_0_i_91 
       (.I0(\slvo[1][hconfig][5] [5]),
        .I1(\slvo[1][hconfig][5] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[1][hconfig][5] [6]),
        .I4(\slvo[1][hconfig][5] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hsel][1]_INST_0_i_91_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \slvi[hsel][2]_INST_0 
       (.I0(p_1_in10_in),
        .I1(hsel1192_out),
        .O(\^slvi[hsel] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFF7F7F7)) 
    \slvi[hsel][2]_INST_0_i_1 
       (.I0(\slvi[hsel][2]_INST_0_i_2_n_0 ),
        .I1(\slvi[hsel][2]_INST_0_i_3_n_0 ),
        .I2(\slvi[hsel][2]_INST_0_i_4_n_0 ),
        .I3(\slvi[hsel][2]_INST_0_i_5_n_0 ),
        .I4(\slvo[2][hconfig][7] [1]),
        .O(p_1_in10_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hsel][2]_INST_0_i_10 
       (.I0(\slvi[hsel][2]_INST_0_i_25_n_0 ),
        .I1(\slvi[hsel][2]_INST_0_i_26_n_0 ),
        .O(hsel2119_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][2]_INST_0_i_11 
       (.CI(slvi),
        .CO({hsel346_out,\slvi[hsel][2]_INST_0_i_11_n_1 ,\slvi[hsel][2]_INST_0_i_11_n_2 ,\slvi[hsel][2]_INST_0_i_11_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][2]_INST_0_i_27_n_0 ,\slvi[hsel][2]_INST_0_i_28_n_0 ,\slvi[hsel][2]_INST_0_i_29_n_0 ,\slvi[hsel][2]_INST_0_i_30_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][2]_INST_0_i_12 
       (.CI(slvi),
        .CO({hsel341_out,\slvi[hsel][2]_INST_0_i_12_n_1 ,\slvi[hsel][2]_INST_0_i_12_n_2 ,\slvi[hsel][2]_INST_0_i_12_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][2]_INST_0_i_31_n_0 ,\slvi[hsel][2]_INST_0_i_32_n_0 ,\slvi[hsel][2]_INST_0_i_33_n_0 ,\slvi[hsel][2]_INST_0_i_34_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hsel][2]_INST_0_i_13 
       (.I0(\slvi[hsel][2]_INST_0_i_35_n_0 ),
        .I1(\slvi[hsel][2]_INST_0_i_36_n_0 ),
        .O(hsel2125_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][2]_INST_0_i_14 
       (.CI(slvi),
        .CO({hsel344_out,\slvi[hsel][2]_INST_0_i_14_n_1 ,\slvi[hsel][2]_INST_0_i_14_n_2 ,\slvi[hsel][2]_INST_0_i_14_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][2]_INST_0_i_37_n_0 ,\slvi[hsel][2]_INST_0_i_38_n_0 ,\slvi[hsel][2]_INST_0_i_39_n_0 ,\slvi[hsel][2]_INST_0_i_40_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][2]_INST_0_i_15 
       (.CI(slvi),
        .CO({hsel342_out,\slvi[hsel][2]_INST_0_i_15_n_1 ,\slvi[hsel][2]_INST_0_i_15_n_2 ,\slvi[hsel][2]_INST_0_i_15_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][2]_INST_0_i_41_n_0 ,\slvi[hsel][2]_INST_0_i_42_n_0 ,\slvi[hsel][2]_INST_0_i_43_n_0 ,\slvi[hsel][2]_INST_0_i_44_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hsel][2]_INST_0_i_16 
       (.I0(\slvi[hsel][2]_INST_0_i_45_n_0 ),
        .I1(\slvi[hsel][2]_INST_0_i_46_n_0 ),
        .O(hsel2128_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][2]_INST_0_i_17 
       (.CI(slvi),
        .CO({hsel343_out,\slvi[hsel][2]_INST_0_i_17_n_1 ,\slvi[hsel][2]_INST_0_i_17_n_2 ,\slvi[hsel][2]_INST_0_i_17_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][2]_INST_0_i_47_n_0 ,\slvi[hsel][2]_INST_0_i_48_n_0 ,\slvi[hsel][2]_INST_0_i_49_n_0 ,\slvi[hsel][2]_INST_0_i_50_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][2]_INST_0_i_18 
       (.CI(slvi),
        .CO({hsel340_out,\slvi[hsel][2]_INST_0_i_18_n_1 ,\slvi[hsel][2]_INST_0_i_18_n_2 ,\slvi[hsel][2]_INST_0_i_18_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][2]_INST_0_i_51_n_0 ,\slvi[hsel][2]_INST_0_i_52_n_0 ,\slvi[hsel][2]_INST_0_i_53_n_0 ,\slvi[hsel][2]_INST_0_i_54_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hsel][2]_INST_0_i_19 
       (.I0(\slvi[hsel][2]_INST_0_i_55_n_0 ),
        .I1(\slvi[hsel][2]_INST_0_i_56_n_0 ),
        .O(hsel2122_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hsel][2]_INST_0_i_2 
       (.I0(\slvo[2][hconfig][5] [1]),
        .I1(\slvi[hsel][2]_INST_0_i_6_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][2]_INST_0_i_20 
       (.CI(slvi),
        .CO({hsel345_out,\slvi[hsel][2]_INST_0_i_20_n_1 ,\slvi[hsel][2]_INST_0_i_20_n_2 ,\slvi[hsel][2]_INST_0_i_20_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][2]_INST_0_i_57_n_0 ,\slvi[hsel][2]_INST_0_i_58_n_0 ,\slvi[hsel][2]_INST_0_i_59_n_0 ,\slvi[hsel][2]_INST_0_i_60_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_21 
       (.I0(\slvo[2][hconfig][7] [13]),
        .I1(\slvo[2][hconfig][7] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hsel][2]_INST_0_i_61_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_22 
       (.I0(\slvo[2][hconfig][7] [10]),
        .I1(\slvo[2][hconfig][7] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hsel][2]_INST_0_i_62_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_23 
       (.I0(\slvo[2][hconfig][7] [7]),
        .I1(\slvo[2][hconfig][7] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hsel][2]_INST_0_i_63_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_24 
       (.I0(\slvo[2][hconfig][7] [4]),
        .I1(\slvo[2][hconfig][7] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hsel][2]_INST_0_i_64_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][2]_INST_0_i_25 
       (.I0(\slvo[2][hconfig][7] [9]),
        .I1(\slvo[2][hconfig][7] [7]),
        .I2(\slvo[2][hconfig][7] [8]),
        .I3(\slvo[2][hconfig][7] [4]),
        .I4(\slvo[2][hconfig][7] [5]),
        .I5(\slvo[2][hconfig][7] [6]),
        .O(\slvi[hsel][2]_INST_0_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][2]_INST_0_i_26 
       (.I0(\slvo[2][hconfig][7] [14]),
        .I1(\slvo[2][hconfig][7] [13]),
        .I2(\slvo[2][hconfig][7] [15]),
        .I3(\slvo[2][hconfig][7] [10]),
        .I4(\slvo[2][hconfig][7] [11]),
        .I5(\slvo[2][hconfig][7] [12]),
        .O(\slvi[hsel][2]_INST_0_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_27 
       (.I0(\slvo[2][hconfig][7] [13]),
        .I1(\slvo[2][hconfig][7] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hsel][2]_INST_0_i_65_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_28 
       (.I0(\slvo[2][hconfig][7] [10]),
        .I1(\slvo[2][hconfig][7] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hsel][2]_INST_0_i_66_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_29 
       (.I0(\slvo[2][hconfig][7] [7]),
        .I1(\slvo[2][hconfig][7] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hsel][2]_INST_0_i_67_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hsel][2]_INST_0_i_3 
       (.I0(\slvo[2][hconfig][4] [1]),
        .I1(\slvi[hsel][2]_INST_0_i_7_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_30 
       (.I0(\slvo[2][hconfig][7] [4]),
        .I1(\slvo[2][hconfig][7] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hsel][2]_INST_0_i_68_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_31 
       (.I0(\slvo[2][hconfig][5] [13]),
        .I1(\slvo[2][hconfig][5] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hsel][2]_INST_0_i_69_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_32 
       (.I0(\slvo[2][hconfig][5] [10]),
        .I1(\slvo[2][hconfig][5] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hsel][2]_INST_0_i_70_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_33 
       (.I0(\slvo[2][hconfig][5] [7]),
        .I1(\slvo[2][hconfig][5] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hsel][2]_INST_0_i_71_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_34 
       (.I0(\slvo[2][hconfig][5] [4]),
        .I1(\slvo[2][hconfig][5] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hsel][2]_INST_0_i_72_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][2]_INST_0_i_35 
       (.I0(\slvo[2][hconfig][5] [9]),
        .I1(\slvo[2][hconfig][5] [7]),
        .I2(\slvo[2][hconfig][5] [8]),
        .I3(\slvo[2][hconfig][5] [4]),
        .I4(\slvo[2][hconfig][5] [5]),
        .I5(\slvo[2][hconfig][5] [6]),
        .O(\slvi[hsel][2]_INST_0_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][2]_INST_0_i_36 
       (.I0(\slvo[2][hconfig][5] [14]),
        .I1(\slvo[2][hconfig][5] [13]),
        .I2(\slvo[2][hconfig][5] [15]),
        .I3(\slvo[2][hconfig][5] [10]),
        .I4(\slvo[2][hconfig][5] [11]),
        .I5(\slvo[2][hconfig][5] [12]),
        .O(\slvi[hsel][2]_INST_0_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_37 
       (.I0(\slvo[2][hconfig][5] [13]),
        .I1(\slvo[2][hconfig][5] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hsel][2]_INST_0_i_73_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_38 
       (.I0(\slvo[2][hconfig][5] [10]),
        .I1(\slvo[2][hconfig][5] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hsel][2]_INST_0_i_74_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_39 
       (.I0(\slvo[2][hconfig][5] [7]),
        .I1(\slvo[2][hconfig][5] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hsel][2]_INST_0_i_75_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \slvi[hsel][2]_INST_0_i_4 
       (.I0(\slvi[hsel][2]_INST_0_i_8_n_0 ),
        .I1(\slvo[2][hconfig][6] [1]),
        .O(\slvi[hsel][2]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_40 
       (.I0(\slvo[2][hconfig][5] [4]),
        .I1(\slvo[2][hconfig][5] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hsel][2]_INST_0_i_76_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_41 
       (.I0(\slvo[2][hconfig][4] [13]),
        .I1(\slvo[2][hconfig][4] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hsel][2]_INST_0_i_77_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_42 
       (.I0(\slvo[2][hconfig][4] [10]),
        .I1(\slvo[2][hconfig][4] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hsel][2]_INST_0_i_78_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_43 
       (.I0(\slvo[2][hconfig][4] [7]),
        .I1(\slvo[2][hconfig][4] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hsel][2]_INST_0_i_79_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_44 
       (.I0(\slvo[2][hconfig][4] [4]),
        .I1(\slvo[2][hconfig][4] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hsel][2]_INST_0_i_80_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][2]_INST_0_i_45 
       (.I0(\slvo[2][hconfig][4] [9]),
        .I1(\slvo[2][hconfig][4] [7]),
        .I2(\slvo[2][hconfig][4] [8]),
        .I3(\slvo[2][hconfig][4] [4]),
        .I4(\slvo[2][hconfig][4] [5]),
        .I5(\slvo[2][hconfig][4] [6]),
        .O(\slvi[hsel][2]_INST_0_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][2]_INST_0_i_46 
       (.I0(\slvo[2][hconfig][4] [14]),
        .I1(\slvo[2][hconfig][4] [13]),
        .I2(\slvo[2][hconfig][4] [15]),
        .I3(\slvo[2][hconfig][4] [10]),
        .I4(\slvo[2][hconfig][4] [11]),
        .I5(\slvo[2][hconfig][4] [12]),
        .O(\slvi[hsel][2]_INST_0_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_47 
       (.I0(\slvo[2][hconfig][4] [13]),
        .I1(\slvo[2][hconfig][4] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hsel][2]_INST_0_i_81_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_48 
       (.I0(\slvo[2][hconfig][4] [10]),
        .I1(\slvo[2][hconfig][4] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hsel][2]_INST_0_i_82_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_49 
       (.I0(\slvo[2][hconfig][4] [7]),
        .I1(\slvo[2][hconfig][4] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hsel][2]_INST_0_i_83_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h80808080F0000000)) 
    \slvi[hsel][2]_INST_0_i_5 
       (.I0(hsel339_out),
        .I1(hsel219_in),
        .I2(hsel2119_in),
        .I3(hsel346_out),
        .I4(hsel330_in),
        .I5(\slvo[2][hconfig][7] [0]),
        .O(\slvi[hsel][2]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_50 
       (.I0(\slvo[2][hconfig][4] [4]),
        .I1(\slvo[2][hconfig][4] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hsel][2]_INST_0_i_84_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_51 
       (.I0(\slvo[2][hconfig][6] [13]),
        .I1(\slvo[2][hconfig][6] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hsel][2]_INST_0_i_85_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_51_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_52 
       (.I0(\slvo[2][hconfig][6] [10]),
        .I1(\slvo[2][hconfig][6] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hsel][2]_INST_0_i_86_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_52_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_53 
       (.I0(\slvo[2][hconfig][6] [7]),
        .I1(\slvo[2][hconfig][6] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hsel][2]_INST_0_i_87_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_53_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_54 
       (.I0(\slvo[2][hconfig][6] [4]),
        .I1(\slvo[2][hconfig][6] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hsel][2]_INST_0_i_88_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_54_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][2]_INST_0_i_55 
       (.I0(\slvo[2][hconfig][6] [9]),
        .I1(\slvo[2][hconfig][6] [7]),
        .I2(\slvo[2][hconfig][6] [8]),
        .I3(\slvo[2][hconfig][6] [4]),
        .I4(\slvo[2][hconfig][6] [5]),
        .I5(\slvo[2][hconfig][6] [6]),
        .O(\slvi[hsel][2]_INST_0_i_55_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][2]_INST_0_i_56 
       (.I0(\slvo[2][hconfig][6] [14]),
        .I1(\slvo[2][hconfig][6] [13]),
        .I2(\slvo[2][hconfig][6] [15]),
        .I3(\slvo[2][hconfig][6] [10]),
        .I4(\slvo[2][hconfig][6] [11]),
        .I5(\slvo[2][hconfig][6] [12]),
        .O(\slvi[hsel][2]_INST_0_i_56_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_57 
       (.I0(\slvo[2][hconfig][6] [13]),
        .I1(\slvo[2][hconfig][6] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hsel][2]_INST_0_i_89_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_57_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_58 
       (.I0(\slvo[2][hconfig][6] [10]),
        .I1(\slvo[2][hconfig][6] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hsel][2]_INST_0_i_90_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_58_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_59 
       (.I0(\slvo[2][hconfig][6] [7]),
        .I1(\slvo[2][hconfig][6] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hsel][2]_INST_0_i_91_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_59_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000808030003000)) 
    \slvi[hsel][2]_INST_0_i_6 
       (.I0(hsel341_out),
        .I1(\slvo[2][hconfig][5] [0]),
        .I2(hsel2125_in),
        .I3(hsel344_out),
        .I4(\slvi[hmbsel][2]_INST_0_i_9_n_0 ),
        .I5(\slvi[hmbsel][2]_INST_0_i_10_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][2]_INST_0_i_60 
       (.I0(\slvo[2][hconfig][6] [4]),
        .I1(\slvo[2][hconfig][6] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hsel][2]_INST_0_i_92_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_60_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_61 
       (.I0(\slvo[2][hconfig][7] [14]),
        .I1(\slvo[2][hconfig][7] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[2][hconfig][7] [15]),
        .I4(\slvo[2][hconfig][7] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hsel][2]_INST_0_i_61_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_62 
       (.I0(\slvo[2][hconfig][7] [11]),
        .I1(\slvo[2][hconfig][7] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[2][hconfig][7] [12]),
        .I4(\slvo[2][hconfig][7] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hsel][2]_INST_0_i_62_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_63 
       (.I0(\slvo[2][hconfig][7] [8]),
        .I1(\slvo[2][hconfig][7] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[2][hconfig][7] [9]),
        .I4(\slvo[2][hconfig][7] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hsel][2]_INST_0_i_63_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_64 
       (.I0(\slvo[2][hconfig][7] [5]),
        .I1(\slvo[2][hconfig][7] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[2][hconfig][7] [6]),
        .I4(\slvo[2][hconfig][7] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hsel][2]_INST_0_i_64_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_65 
       (.I0(\slvo[2][hconfig][7] [14]),
        .I1(\slvo[2][hconfig][7] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[2][hconfig][7] [15]),
        .I4(\slvo[2][hconfig][7] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hsel][2]_INST_0_i_65_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_66 
       (.I0(\slvo[2][hconfig][7] [11]),
        .I1(\slvo[2][hconfig][7] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[2][hconfig][7] [12]),
        .I4(\slvo[2][hconfig][7] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hsel][2]_INST_0_i_66_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_67 
       (.I0(\slvo[2][hconfig][7] [8]),
        .I1(\slvo[2][hconfig][7] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[2][hconfig][7] [9]),
        .I4(\slvo[2][hconfig][7] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hsel][2]_INST_0_i_67_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_68 
       (.I0(\slvo[2][hconfig][7] [5]),
        .I1(\slvo[2][hconfig][7] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[2][hconfig][7] [6]),
        .I4(\slvo[2][hconfig][7] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hsel][2]_INST_0_i_68_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_69 
       (.I0(\slvo[2][hconfig][5] [14]),
        .I1(\slvo[2][hconfig][5] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[2][hconfig][5] [15]),
        .I4(\slvo[2][hconfig][5] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hsel][2]_INST_0_i_69_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000808030003000)) 
    \slvi[hsel][2]_INST_0_i_7 
       (.I0(hsel342_out),
        .I1(\slvo[2][hconfig][4] [0]),
        .I2(hsel2128_in),
        .I3(hsel343_out),
        .I4(\slvi[hmbsel][2]_INST_0_i_9_n_0 ),
        .I5(\slvi[hmbsel][2]_INST_0_i_10_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_70 
       (.I0(\slvo[2][hconfig][5] [11]),
        .I1(\slvo[2][hconfig][5] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[2][hconfig][5] [12]),
        .I4(\slvo[2][hconfig][5] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hsel][2]_INST_0_i_70_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_71 
       (.I0(\slvo[2][hconfig][5] [8]),
        .I1(\slvo[2][hconfig][5] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[2][hconfig][5] [9]),
        .I4(\slvo[2][hconfig][5] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hsel][2]_INST_0_i_71_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_72 
       (.I0(\slvo[2][hconfig][5] [5]),
        .I1(\slvo[2][hconfig][5] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[2][hconfig][5] [6]),
        .I4(\slvo[2][hconfig][5] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hsel][2]_INST_0_i_72_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_73 
       (.I0(\slvo[2][hconfig][5] [14]),
        .I1(\slvo[2][hconfig][5] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[2][hconfig][5] [15]),
        .I4(\slvo[2][hconfig][5] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hsel][2]_INST_0_i_73_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_74 
       (.I0(\slvo[2][hconfig][5] [11]),
        .I1(\slvo[2][hconfig][5] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[2][hconfig][5] [12]),
        .I4(\slvo[2][hconfig][5] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hsel][2]_INST_0_i_74_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_75 
       (.I0(\slvo[2][hconfig][5] [8]),
        .I1(\slvo[2][hconfig][5] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[2][hconfig][5] [9]),
        .I4(\slvo[2][hconfig][5] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hsel][2]_INST_0_i_75_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_76 
       (.I0(\slvo[2][hconfig][5] [5]),
        .I1(\slvo[2][hconfig][5] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[2][hconfig][5] [6]),
        .I4(\slvo[2][hconfig][5] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hsel][2]_INST_0_i_76_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_77 
       (.I0(\slvo[2][hconfig][4] [14]),
        .I1(\slvo[2][hconfig][4] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[2][hconfig][4] [15]),
        .I4(\slvo[2][hconfig][4] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hsel][2]_INST_0_i_77_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_78 
       (.I0(\slvo[2][hconfig][4] [11]),
        .I1(\slvo[2][hconfig][4] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[2][hconfig][4] [12]),
        .I4(\slvo[2][hconfig][4] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hsel][2]_INST_0_i_78_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_79 
       (.I0(\slvo[2][hconfig][4] [8]),
        .I1(\slvo[2][hconfig][4] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[2][hconfig][4] [9]),
        .I4(\slvo[2][hconfig][4] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hsel][2]_INST_0_i_79_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000808030003000)) 
    \slvi[hsel][2]_INST_0_i_8 
       (.I0(hsel340_out),
        .I1(\slvo[2][hconfig][6] [0]),
        .I2(hsel2122_in),
        .I3(hsel345_out),
        .I4(\slvi[hmbsel][2]_INST_0_i_9_n_0 ),
        .I5(\slvi[hmbsel][2]_INST_0_i_10_n_0 ),
        .O(\slvi[hsel][2]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_80 
       (.I0(\slvo[2][hconfig][4] [5]),
        .I1(\slvo[2][hconfig][4] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[2][hconfig][4] [6]),
        .I4(\slvo[2][hconfig][4] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hsel][2]_INST_0_i_80_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_81 
       (.I0(\slvo[2][hconfig][4] [14]),
        .I1(\slvo[2][hconfig][4] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[2][hconfig][4] [15]),
        .I4(\slvo[2][hconfig][4] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hsel][2]_INST_0_i_81_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_82 
       (.I0(\slvo[2][hconfig][4] [11]),
        .I1(\slvo[2][hconfig][4] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[2][hconfig][4] [12]),
        .I4(\slvo[2][hconfig][4] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hsel][2]_INST_0_i_82_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_83 
       (.I0(\slvo[2][hconfig][4] [8]),
        .I1(\slvo[2][hconfig][4] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[2][hconfig][4] [9]),
        .I4(\slvo[2][hconfig][4] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hsel][2]_INST_0_i_83_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_84 
       (.I0(\slvo[2][hconfig][4] [5]),
        .I1(\slvo[2][hconfig][4] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[2][hconfig][4] [6]),
        .I4(\slvo[2][hconfig][4] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hsel][2]_INST_0_i_84_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_85 
       (.I0(\slvo[2][hconfig][6] [14]),
        .I1(\slvo[2][hconfig][6] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[2][hconfig][6] [15]),
        .I4(\slvo[2][hconfig][6] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hsel][2]_INST_0_i_85_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_86 
       (.I0(\slvo[2][hconfig][6] [11]),
        .I1(\slvo[2][hconfig][6] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[2][hconfig][6] [12]),
        .I4(\slvo[2][hconfig][6] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hsel][2]_INST_0_i_86_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_87 
       (.I0(\slvo[2][hconfig][6] [8]),
        .I1(\slvo[2][hconfig][6] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[2][hconfig][6] [9]),
        .I4(\slvo[2][hconfig][6] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hsel][2]_INST_0_i_87_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_88 
       (.I0(\slvo[2][hconfig][6] [5]),
        .I1(\slvo[2][hconfig][6] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[2][hconfig][6] [6]),
        .I4(\slvo[2][hconfig][6] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hsel][2]_INST_0_i_88_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_89 
       (.I0(\slvo[2][hconfig][6] [14]),
        .I1(\slvo[2][hconfig][6] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[2][hconfig][6] [15]),
        .I4(\slvo[2][hconfig][6] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hsel][2]_INST_0_i_89_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][2]_INST_0_i_9 
       (.CI(slvi),
        .CO({hsel339_out,\slvi[hsel][2]_INST_0_i_9_n_1 ,\slvi[hsel][2]_INST_0_i_9_n_2 ,\slvi[hsel][2]_INST_0_i_9_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][2]_INST_0_i_21_n_0 ,\slvi[hsel][2]_INST_0_i_22_n_0 ,\slvi[hsel][2]_INST_0_i_23_n_0 ,\slvi[hsel][2]_INST_0_i_24_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_90 
       (.I0(\slvo[2][hconfig][6] [11]),
        .I1(\slvo[2][hconfig][6] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[2][hconfig][6] [12]),
        .I4(\slvo[2][hconfig][6] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hsel][2]_INST_0_i_90_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_91 
       (.I0(\slvo[2][hconfig][6] [8]),
        .I1(\slvo[2][hconfig][6] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[2][hconfig][6] [9]),
        .I4(\slvo[2][hconfig][6] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hsel][2]_INST_0_i_91_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][2]_INST_0_i_92 
       (.I0(\slvo[2][hconfig][6] [5]),
        .I1(\slvo[2][hconfig][6] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[2][hconfig][6] [6]),
        .I4(\slvo[2][hconfig][6] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hsel][2]_INST_0_i_92_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \slvi[hsel][3]_INST_0 
       (.I0(p_0_in5_in),
        .I1(hsel1192_out),
        .O(\^slvi[hsel] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFF7F7F7)) 
    \slvi[hsel][3]_INST_0_i_1 
       (.I0(\slvi[hmbsel][1]_INST_0_i_4_n_0 ),
        .I1(\slvi[hmbsel][0]_INST_0_i_4_n_0 ),
        .I2(\slvi[hsel][3]_INST_0_i_2_n_0 ),
        .I3(\slvi[hsel][3]_INST_0_i_3_n_0 ),
        .I4(\slvo[3][hconfig][7] [1]),
        .O(p_0_in5_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][3]_INST_0_i_10 
       (.CI(slvi),
        .CO({hsel337_out,\slvi[hsel][3]_INST_0_i_10_n_1 ,\slvi[hsel][3]_INST_0_i_10_n_2 ,\slvi[hsel][3]_INST_0_i_10_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][3]_INST_0_i_27_n_0 ,\slvi[hsel][3]_INST_0_i_28_n_0 ,\slvi[hsel][3]_INST_0_i_29_n_0 ,\slvi[hsel][3]_INST_0_i_30_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][3]_INST_0_i_11 
       (.I0(\slvo[3][hconfig][7] [13]),
        .I1(\slvo[3][hconfig][7] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hsel][3]_INST_0_i_31_n_0 ),
        .O(\slvi[hsel][3]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][3]_INST_0_i_12 
       (.I0(\slvo[3][hconfig][7] [10]),
        .I1(\slvo[3][hconfig][7] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hsel][3]_INST_0_i_32_n_0 ),
        .O(\slvi[hsel][3]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][3]_INST_0_i_13 
       (.I0(\slvo[3][hconfig][7] [7]),
        .I1(\slvo[3][hconfig][7] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hsel][3]_INST_0_i_33_n_0 ),
        .O(\slvi[hsel][3]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][3]_INST_0_i_14 
       (.I0(\slvo[3][hconfig][7] [4]),
        .I1(\slvo[3][hconfig][7] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hsel][3]_INST_0_i_34_n_0 ),
        .O(\slvi[hsel][3]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][3]_INST_0_i_15 
       (.I0(\slvo[3][hconfig][7] [9]),
        .I1(\slvo[3][hconfig][7] [7]),
        .I2(\slvo[3][hconfig][7] [8]),
        .I3(\slvo[3][hconfig][7] [4]),
        .I4(\slvo[3][hconfig][7] [5]),
        .I5(\slvo[3][hconfig][7] [6]),
        .O(\slvi[hsel][3]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][3]_INST_0_i_16 
       (.I0(\slvo[3][hconfig][7] [14]),
        .I1(\slvo[3][hconfig][7] [13]),
        .I2(\slvo[3][hconfig][7] [15]),
        .I3(\slvo[3][hconfig][7] [10]),
        .I4(\slvo[3][hconfig][7] [11]),
        .I5(\slvo[3][hconfig][7] [12]),
        .O(\slvi[hsel][3]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][3]_INST_0_i_17 
       (.I0(\slvo[3][hconfig][7] [13]),
        .I1(\slvo[3][hconfig][7] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hsel][3]_INST_0_i_35_n_0 ),
        .O(\slvi[hsel][3]_INST_0_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][3]_INST_0_i_18 
       (.I0(\slvo[3][hconfig][7] [10]),
        .I1(\slvo[3][hconfig][7] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hsel][3]_INST_0_i_36_n_0 ),
        .O(\slvi[hsel][3]_INST_0_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][3]_INST_0_i_19 
       (.I0(\slvo[3][hconfig][7] [7]),
        .I1(\slvo[3][hconfig][7] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hsel][3]_INST_0_i_37_n_0 ),
        .O(\slvi[hsel][3]_INST_0_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \slvi[hsel][3]_INST_0_i_2 
       (.I0(\slvi[hsel][3]_INST_0_i_4_n_0 ),
        .I1(\slvo[3][hconfig][6] [1]),
        .O(\slvi[hsel][3]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][3]_INST_0_i_20 
       (.I0(\slvo[3][hconfig][7] [4]),
        .I1(\slvo[3][hconfig][7] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hsel][3]_INST_0_i_38_n_0 ),
        .O(\slvi[hsel][3]_INST_0_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][3]_INST_0_i_21 
       (.I0(\slvo[3][hconfig][6] [13]),
        .I1(\slvo[3][hconfig][6] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hsel][3]_INST_0_i_39_n_0 ),
        .O(\slvi[hsel][3]_INST_0_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][3]_INST_0_i_22 
       (.I0(\slvo[3][hconfig][6] [10]),
        .I1(\slvo[3][hconfig][6] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hsel][3]_INST_0_i_40_n_0 ),
        .O(\slvi[hsel][3]_INST_0_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][3]_INST_0_i_23 
       (.I0(\slvo[3][hconfig][6] [7]),
        .I1(\slvo[3][hconfig][6] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hsel][3]_INST_0_i_41_n_0 ),
        .O(\slvi[hsel][3]_INST_0_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][3]_INST_0_i_24 
       (.I0(\slvo[3][hconfig][6] [4]),
        .I1(\slvo[3][hconfig][6] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hsel][3]_INST_0_i_42_n_0 ),
        .O(\slvi[hsel][3]_INST_0_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][3]_INST_0_i_25 
       (.I0(\slvo[3][hconfig][6] [9]),
        .I1(\slvo[3][hconfig][6] [7]),
        .I2(\slvo[3][hconfig][6] [8]),
        .I3(\slvo[3][hconfig][6] [4]),
        .I4(\slvo[3][hconfig][6] [5]),
        .I5(\slvo[3][hconfig][6] [6]),
        .O(\slvi[hsel][3]_INST_0_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][3]_INST_0_i_26 
       (.I0(\slvo[3][hconfig][6] [14]),
        .I1(\slvo[3][hconfig][6] [13]),
        .I2(\slvo[3][hconfig][6] [15]),
        .I3(\slvo[3][hconfig][6] [10]),
        .I4(\slvo[3][hconfig][6] [11]),
        .I5(\slvo[3][hconfig][6] [12]),
        .O(\slvi[hsel][3]_INST_0_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][3]_INST_0_i_27 
       (.I0(\slvo[3][hconfig][6] [13]),
        .I1(\slvo[3][hconfig][6] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hsel][3]_INST_0_i_43_n_0 ),
        .O(\slvi[hsel][3]_INST_0_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][3]_INST_0_i_28 
       (.I0(\slvo[3][hconfig][6] [10]),
        .I1(\slvo[3][hconfig][6] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hsel][3]_INST_0_i_44_n_0 ),
        .O(\slvi[hsel][3]_INST_0_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][3]_INST_0_i_29 
       (.I0(\slvo[3][hconfig][6] [7]),
        .I1(\slvo[3][hconfig][6] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hsel][3]_INST_0_i_45_n_0 ),
        .O(\slvi[hsel][3]_INST_0_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h80808080F0000000)) 
    \slvi[hsel][3]_INST_0_i_3 
       (.I0(hsel331_out),
        .I1(hsel219_in),
        .I2(hsel299_in),
        .I3(hsel338_out),
        .I4(hsel330_in),
        .I5(\slvo[3][hconfig][7] [0]),
        .O(\slvi[hsel][3]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][3]_INST_0_i_30 
       (.I0(\slvo[3][hconfig][6] [4]),
        .I1(\slvo[3][hconfig][6] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hsel][3]_INST_0_i_46_n_0 ),
        .O(\slvi[hsel][3]_INST_0_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][3]_INST_0_i_31 
       (.I0(\slvo[3][hconfig][7] [14]),
        .I1(\slvo[3][hconfig][7] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[3][hconfig][7] [15]),
        .I4(\slvo[3][hconfig][7] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hsel][3]_INST_0_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][3]_INST_0_i_32 
       (.I0(\slvo[3][hconfig][7] [11]),
        .I1(\slvo[3][hconfig][7] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[3][hconfig][7] [12]),
        .I4(\slvo[3][hconfig][7] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hsel][3]_INST_0_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][3]_INST_0_i_33 
       (.I0(\slvo[3][hconfig][7] [8]),
        .I1(\slvo[3][hconfig][7] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[3][hconfig][7] [9]),
        .I4(\slvo[3][hconfig][7] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hsel][3]_INST_0_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][3]_INST_0_i_34 
       (.I0(\slvo[3][hconfig][7] [5]),
        .I1(\slvo[3][hconfig][7] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[3][hconfig][7] [6]),
        .I4(\slvo[3][hconfig][7] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hsel][3]_INST_0_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][3]_INST_0_i_35 
       (.I0(\slvo[3][hconfig][7] [14]),
        .I1(\slvo[3][hconfig][7] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[3][hconfig][7] [15]),
        .I4(\slvo[3][hconfig][7] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hsel][3]_INST_0_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][3]_INST_0_i_36 
       (.I0(\slvo[3][hconfig][7] [11]),
        .I1(\slvo[3][hconfig][7] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[3][hconfig][7] [12]),
        .I4(\slvo[3][hconfig][7] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hsel][3]_INST_0_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][3]_INST_0_i_37 
       (.I0(\slvo[3][hconfig][7] [8]),
        .I1(\slvo[3][hconfig][7] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[3][hconfig][7] [9]),
        .I4(\slvo[3][hconfig][7] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hsel][3]_INST_0_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][3]_INST_0_i_38 
       (.I0(\slvo[3][hconfig][7] [5]),
        .I1(\slvo[3][hconfig][7] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[3][hconfig][7] [6]),
        .I4(\slvo[3][hconfig][7] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hsel][3]_INST_0_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][3]_INST_0_i_39 
       (.I0(\slvo[3][hconfig][6] [14]),
        .I1(\slvo[3][hconfig][6] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[3][hconfig][6] [15]),
        .I4(\slvo[3][hconfig][6] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hsel][3]_INST_0_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000808030003000)) 
    \slvi[hsel][3]_INST_0_i_4 
       (.I0(hsel332_out),
        .I1(\slvo[3][hconfig][6] [0]),
        .I2(hsel2102_in),
        .I3(hsel337_out),
        .I4(\slvi[hmbsel][2]_INST_0_i_9_n_0 ),
        .I5(\slvi[hmbsel][2]_INST_0_i_10_n_0 ),
        .O(\slvi[hsel][3]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][3]_INST_0_i_40 
       (.I0(\slvo[3][hconfig][6] [11]),
        .I1(\slvo[3][hconfig][6] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[3][hconfig][6] [12]),
        .I4(\slvo[3][hconfig][6] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hsel][3]_INST_0_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][3]_INST_0_i_41 
       (.I0(\slvo[3][hconfig][6] [8]),
        .I1(\slvo[3][hconfig][6] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[3][hconfig][6] [9]),
        .I4(\slvo[3][hconfig][6] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hsel][3]_INST_0_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][3]_INST_0_i_42 
       (.I0(\slvo[3][hconfig][6] [5]),
        .I1(\slvo[3][hconfig][6] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[3][hconfig][6] [6]),
        .I4(\slvo[3][hconfig][6] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hsel][3]_INST_0_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][3]_INST_0_i_43 
       (.I0(\slvo[3][hconfig][6] [14]),
        .I1(\slvo[3][hconfig][6] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[3][hconfig][6] [15]),
        .I4(\slvo[3][hconfig][6] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hsel][3]_INST_0_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][3]_INST_0_i_44 
       (.I0(\slvo[3][hconfig][6] [11]),
        .I1(\slvo[3][hconfig][6] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[3][hconfig][6] [12]),
        .I4(\slvo[3][hconfig][6] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hsel][3]_INST_0_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][3]_INST_0_i_45 
       (.I0(\slvo[3][hconfig][6] [8]),
        .I1(\slvo[3][hconfig][6] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[3][hconfig][6] [9]),
        .I4(\slvo[3][hconfig][6] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hsel][3]_INST_0_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][3]_INST_0_i_46 
       (.I0(\slvo[3][hconfig][6] [5]),
        .I1(\slvo[3][hconfig][6] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[3][hconfig][6] [6]),
        .I4(\slvo[3][hconfig][6] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hsel][3]_INST_0_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][3]_INST_0_i_5 
       (.CI(slvi),
        .CO({hsel331_out,\slvi[hsel][3]_INST_0_i_5_n_1 ,\slvi[hsel][3]_INST_0_i_5_n_2 ,\slvi[hsel][3]_INST_0_i_5_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][3]_INST_0_i_11_n_0 ,\slvi[hsel][3]_INST_0_i_12_n_0 ,\slvi[hsel][3]_INST_0_i_13_n_0 ,\slvi[hsel][3]_INST_0_i_14_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hsel][3]_INST_0_i_6 
       (.I0(\slvi[hsel][3]_INST_0_i_15_n_0 ),
        .I1(\slvi[hsel][3]_INST_0_i_16_n_0 ),
        .O(hsel299_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][3]_INST_0_i_7 
       (.CI(slvi),
        .CO({hsel338_out,\slvi[hsel][3]_INST_0_i_7_n_1 ,\slvi[hsel][3]_INST_0_i_7_n_2 ,\slvi[hsel][3]_INST_0_i_7_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][3]_INST_0_i_17_n_0 ,\slvi[hsel][3]_INST_0_i_18_n_0 ,\slvi[hsel][3]_INST_0_i_19_n_0 ,\slvi[hsel][3]_INST_0_i_20_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][3]_INST_0_i_8 
       (.CI(slvi),
        .CO({hsel332_out,\slvi[hsel][3]_INST_0_i_8_n_1 ,\slvi[hsel][3]_INST_0_i_8_n_2 ,\slvi[hsel][3]_INST_0_i_8_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][3]_INST_0_i_21_n_0 ,\slvi[hsel][3]_INST_0_i_22_n_0 ,\slvi[hsel][3]_INST_0_i_23_n_0 ,\slvi[hsel][3]_INST_0_i_24_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hsel][3]_INST_0_i_9 
       (.I0(\slvi[hsel][3]_INST_0_i_25_n_0 ),
        .I1(\slvi[hsel][3]_INST_0_i_26_n_0 ),
        .O(hsel2102_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \slvi[hsel][4]_INST_0 
       (.I0(p_1_in13_in),
        .I1(hsel1192_out),
        .O(\^slvi[hsel] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFF7F7F7)) 
    \slvi[hsel][4]_INST_0_i_1 
       (.I0(\slvi[hmbsel][1]_INST_0_i_2_n_0 ),
        .I1(\slvi[hmbsel][0]_INST_0_i_2_n_0 ),
        .I2(\slvi[hmbsel][2]_INST_0_i_3_n_0 ),
        .I3(\slvi[hsel][4]_INST_0_i_2_n_0 ),
        .I4(\slvo[4][hconfig][7] [1]),
        .O(p_1_in13_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][4]_INST_0_i_10 
       (.I0(\slvo[4][hconfig][7] [9]),
        .I1(\slvo[4][hconfig][7] [7]),
        .I2(\slvo[4][hconfig][7] [8]),
        .I3(\slvo[4][hconfig][7] [4]),
        .I4(\slvo[4][hconfig][7] [5]),
        .I5(\slvo[4][hconfig][7] [6]),
        .O(\slvi[hsel][4]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][4]_INST_0_i_11 
       (.I0(\slvo[4][hconfig][7] [14]),
        .I1(\slvo[4][hconfig][7] [13]),
        .I2(\slvo[4][hconfig][7] [15]),
        .I3(\slvo[4][hconfig][7] [10]),
        .I4(\slvo[4][hconfig][7] [11]),
        .I5(\slvo[4][hconfig][7] [12]),
        .O(\slvi[hsel][4]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][4]_INST_0_i_12 
       (.I0(\slvo[4][hconfig][7] [13]),
        .I1(\slvo[4][hconfig][7] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hsel][4]_INST_0_i_20_n_0 ),
        .O(\slvi[hsel][4]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][4]_INST_0_i_13 
       (.I0(\slvo[4][hconfig][7] [10]),
        .I1(\slvo[4][hconfig][7] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hsel][4]_INST_0_i_21_n_0 ),
        .O(\slvi[hsel][4]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][4]_INST_0_i_14 
       (.I0(\slvo[4][hconfig][7] [7]),
        .I1(\slvo[4][hconfig][7] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hsel][4]_INST_0_i_22_n_0 ),
        .O(\slvi[hsel][4]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][4]_INST_0_i_15 
       (.I0(\slvo[4][hconfig][7] [4]),
        .I1(\slvo[4][hconfig][7] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hsel][4]_INST_0_i_23_n_0 ),
        .O(\slvi[hsel][4]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][4]_INST_0_i_16 
       (.I0(\slvo[4][hconfig][7] [14]),
        .I1(\slvo[4][hconfig][7] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[4][hconfig][7] [15]),
        .I4(\slvo[4][hconfig][7] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hsel][4]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][4]_INST_0_i_17 
       (.I0(\slvo[4][hconfig][7] [11]),
        .I1(\slvo[4][hconfig][7] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[4][hconfig][7] [12]),
        .I4(\slvo[4][hconfig][7] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hsel][4]_INST_0_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][4]_INST_0_i_18 
       (.I0(\slvo[4][hconfig][7] [8]),
        .I1(\slvo[4][hconfig][7] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[4][hconfig][7] [9]),
        .I4(\slvo[4][hconfig][7] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hsel][4]_INST_0_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][4]_INST_0_i_19 
       (.I0(\slvo[4][hconfig][7] [5]),
        .I1(\slvo[4][hconfig][7] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[4][hconfig][7] [6]),
        .I4(\slvo[4][hconfig][7] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hsel][4]_INST_0_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h80808080F0000000)) 
    \slvi[hsel][4]_INST_0_i_2 
       (.I0(hsel323_out),
        .I1(hsel219_in),
        .I2(hsel279_in),
        .I3(hsel330_out),
        .I4(hsel330_in),
        .I5(\slvo[4][hconfig][7] [0]),
        .O(\slvi[hsel][4]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][4]_INST_0_i_20 
       (.I0(\slvo[4][hconfig][7] [14]),
        .I1(\slvo[4][hconfig][7] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[4][hconfig][7] [15]),
        .I4(\slvo[4][hconfig][7] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hsel][4]_INST_0_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][4]_INST_0_i_21 
       (.I0(\slvo[4][hconfig][7] [11]),
        .I1(\slvo[4][hconfig][7] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[4][hconfig][7] [12]),
        .I4(\slvo[4][hconfig][7] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hsel][4]_INST_0_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][4]_INST_0_i_22 
       (.I0(\slvo[4][hconfig][7] [8]),
        .I1(\slvo[4][hconfig][7] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[4][hconfig][7] [9]),
        .I4(\slvo[4][hconfig][7] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hsel][4]_INST_0_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][4]_INST_0_i_23 
       (.I0(\slvo[4][hconfig][7] [5]),
        .I1(\slvo[4][hconfig][7] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[4][hconfig][7] [6]),
        .I4(\slvo[4][hconfig][7] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hsel][4]_INST_0_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][4]_INST_0_i_3 
       (.CI(slvi),
        .CO({hsel323_out,\slvi[hsel][4]_INST_0_i_3_n_1 ,\slvi[hsel][4]_INST_0_i_3_n_2 ,\slvi[hsel][4]_INST_0_i_3_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][4]_INST_0_i_6_n_0 ,\slvi[hsel][4]_INST_0_i_7_n_0 ,\slvi[hsel][4]_INST_0_i_8_n_0 ,\slvi[hsel][4]_INST_0_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hsel][4]_INST_0_i_4 
       (.I0(\slvi[hsel][4]_INST_0_i_10_n_0 ),
        .I1(\slvi[hsel][4]_INST_0_i_11_n_0 ),
        .O(hsel279_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][4]_INST_0_i_5 
       (.CI(slvi),
        .CO({hsel330_out,\slvi[hsel][4]_INST_0_i_5_n_1 ,\slvi[hsel][4]_INST_0_i_5_n_2 ,\slvi[hsel][4]_INST_0_i_5_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][4]_INST_0_i_12_n_0 ,\slvi[hsel][4]_INST_0_i_13_n_0 ,\slvi[hsel][4]_INST_0_i_14_n_0 ,\slvi[hsel][4]_INST_0_i_15_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][4]_INST_0_i_6 
       (.I0(\slvo[4][hconfig][7] [13]),
        .I1(\slvo[4][hconfig][7] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hsel][4]_INST_0_i_16_n_0 ),
        .O(\slvi[hsel][4]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][4]_INST_0_i_7 
       (.I0(\slvo[4][hconfig][7] [10]),
        .I1(\slvo[4][hconfig][7] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hsel][4]_INST_0_i_17_n_0 ),
        .O(\slvi[hsel][4]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][4]_INST_0_i_8 
       (.I0(\slvo[4][hconfig][7] [7]),
        .I1(\slvo[4][hconfig][7] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hsel][4]_INST_0_i_18_n_0 ),
        .O(\slvi[hsel][4]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][4]_INST_0_i_9 
       (.I0(\slvo[4][hconfig][7] [4]),
        .I1(\slvo[4][hconfig][7] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hsel][4]_INST_0_i_19_n_0 ),
        .O(\slvi[hsel][4]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \slvi[hsel][5]_INST_0 
       (.I0(p_2_in),
        .I1(hsel1192_out),
        .O(\^slvi[hsel] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFF7F7F7)) 
    \slvi[hsel][5]_INST_0_i_1 
       (.I0(\slvi[hmbsel][1]_INST_0_i_5_n_0 ),
        .I1(\slvi[hmbsel][0]_INST_0_i_5_n_0 ),
        .I2(\slvi[hmbsel][2]_INST_0_i_5_n_0 ),
        .I3(\slvi[hsel][5]_INST_0_i_2_n_0 ),
        .I4(\slvo[5][hconfig][7] [1]),
        .O(p_2_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h80808080F0000000)) 
    \slvi[hsel][5]_INST_0_i_2 
       (.I0(hsel315_out),
        .I1(hsel219_in),
        .I2(hsel259_in),
        .I3(hsel322_out),
        .I4(hsel330_in),
        .I5(\slvo[5][hconfig][7] [0]),
        .O(\slvi[hsel][5]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \slvi[hsel][6]_INST_0 
       (.I0(p_2_in7_in),
        .I1(hsel1192_out),
        .O(\^slvi[hsel] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFF7F7F7)) 
    \slvi[hsel][6]_INST_0_i_1 
       (.I0(\slvi[hmbsel][1]_INST_0_i_1_n_0 ),
        .I1(\slvi[hmbsel][0]_INST_0_i_1_n_0 ),
        .I2(\slvi[hmbsel][2]_INST_0_i_2_n_0 ),
        .I3(\slvi[hsel][6]_INST_0_i_2_n_0 ),
        .I4(\slvo[6][hconfig][7] [1]),
        .O(p_2_in7_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h80808080F0000000)) 
    \slvi[hsel][6]_INST_0_i_2 
       (.I0(hsel37_out),
        .I1(hsel219_in),
        .I2(hsel239_in),
        .I3(hsel314_out),
        .I4(hsel330_in),
        .I5(\slvo[6][hconfig][7] [0]),
        .O(\slvi[hsel][6]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \slvi[hsel][7]_INST_0 
       (.I0(\slvi[hsel][7]_INST_0_i_1_n_0 ),
        .I1(hsel1192_out),
        .O(\^slvi[hsel] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h8FFFFFFF)) 
    \slvi[hsel][7]_INST_0_i_1 
       (.I0(\slvo[7][hconfig][6] [1]),
        .I1(\slvi[hmbsel][2]_INST_0_i_1_n_0 ),
        .I2(\slvi[hsel][7]_INST_0_i_2_n_0 ),
        .I3(\slvi[hmbsel][0]_INST_0_i_6_n_0 ),
        .I4(\slvi[hmbsel][1]_INST_0_i_6_n_0 ),
        .O(\slvi[hsel][7]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][7]_INST_0_i_10 
       (.I0(\slvo[7][hconfig][7] [4]),
        .I1(\slvo[7][hconfig][7] [20]),
        .I2(\slvi[haddr] [8]),
        .I3(\slvi[hsel][7]_INST_0_i_20_n_0 ),
        .O(\slvi[hsel][7]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][7]_INST_0_i_11 
       (.I0(\slvo[7][hconfig][7] [9]),
        .I1(\slvo[7][hconfig][7] [7]),
        .I2(\slvo[7][hconfig][7] [8]),
        .I3(\slvo[7][hconfig][7] [4]),
        .I4(\slvo[7][hconfig][7] [5]),
        .I5(\slvo[7][hconfig][7] [6]),
        .O(\slvi[hsel][7]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \slvi[hsel][7]_INST_0_i_12 
       (.I0(\slvo[7][hconfig][7] [14]),
        .I1(\slvo[7][hconfig][7] [13]),
        .I2(\slvo[7][hconfig][7] [15]),
        .I3(\slvo[7][hconfig][7] [10]),
        .I4(\slvo[7][hconfig][7] [11]),
        .I5(\slvo[7][hconfig][7] [12]),
        .O(\slvi[hsel][7]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][7]_INST_0_i_13 
       (.I0(\slvo[7][hconfig][7] [13]),
        .I1(\slvo[7][hconfig][7] [29]),
        .I2(\slvi[haddr] [29]),
        .I3(\slvi[hsel][7]_INST_0_i_21_n_0 ),
        .O(\slvi[hsel][7]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][7]_INST_0_i_14 
       (.I0(\slvo[7][hconfig][7] [10]),
        .I1(\slvo[7][hconfig][7] [26]),
        .I2(\slvi[haddr] [26]),
        .I3(\slvi[hsel][7]_INST_0_i_22_n_0 ),
        .O(\slvi[hsel][7]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][7]_INST_0_i_15 
       (.I0(\slvo[7][hconfig][7] [7]),
        .I1(\slvo[7][hconfig][7] [23]),
        .I2(\slvi[haddr] [23]),
        .I3(\slvi[hsel][7]_INST_0_i_23_n_0 ),
        .O(\slvi[hsel][7]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][7]_INST_0_i_16 
       (.I0(\slvo[7][hconfig][7] [4]),
        .I1(\slvo[7][hconfig][7] [20]),
        .I2(\slvi[haddr] [20]),
        .I3(\slvi[hsel][7]_INST_0_i_24_n_0 ),
        .O(\slvi[hsel][7]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][7]_INST_0_i_17 
       (.I0(\slvo[7][hconfig][7] [14]),
        .I1(\slvo[7][hconfig][7] [30]),
        .I2(\slvi[haddr] [18]),
        .I3(\slvo[7][hconfig][7] [15]),
        .I4(\slvo[7][hconfig][7] [31]),
        .I5(\slvi[haddr] [19]),
        .O(\slvi[hsel][7]_INST_0_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][7]_INST_0_i_18 
       (.I0(\slvo[7][hconfig][7] [11]),
        .I1(\slvo[7][hconfig][7] [27]),
        .I2(\slvi[haddr] [15]),
        .I3(\slvo[7][hconfig][7] [12]),
        .I4(\slvo[7][hconfig][7] [28]),
        .I5(\slvi[haddr] [16]),
        .O(\slvi[hsel][7]_INST_0_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][7]_INST_0_i_19 
       (.I0(\slvo[7][hconfig][7] [8]),
        .I1(\slvo[7][hconfig][7] [24]),
        .I2(\slvi[haddr] [12]),
        .I3(\slvo[7][hconfig][7] [9]),
        .I4(\slvo[7][hconfig][7] [25]),
        .I5(\slvi[haddr] [13]),
        .O(\slvi[hsel][7]_INST_0_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hsel][7]_INST_0_i_2 
       (.I0(\slvo[7][hconfig][7] [1]),
        .I1(\slvi[hsel][7]_INST_0_i_3_n_0 ),
        .O(\slvi[hsel][7]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][7]_INST_0_i_20 
       (.I0(\slvo[7][hconfig][7] [5]),
        .I1(\slvo[7][hconfig][7] [21]),
        .I2(\slvi[haddr] [9]),
        .I3(\slvo[7][hconfig][7] [6]),
        .I4(\slvo[7][hconfig][7] [22]),
        .I5(\slvi[haddr] [10]),
        .O(\slvi[hsel][7]_INST_0_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][7]_INST_0_i_21 
       (.I0(\slvo[7][hconfig][7] [14]),
        .I1(\slvo[7][hconfig][7] [30]),
        .I2(\slvi[haddr] [30]),
        .I3(\slvo[7][hconfig][7] [15]),
        .I4(\slvo[7][hconfig][7] [31]),
        .I5(\slvi[haddr] [31]),
        .O(\slvi[hsel][7]_INST_0_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][7]_INST_0_i_22 
       (.I0(\slvo[7][hconfig][7] [11]),
        .I1(\slvo[7][hconfig][7] [27]),
        .I2(\slvi[haddr] [27]),
        .I3(\slvo[7][hconfig][7] [12]),
        .I4(\slvo[7][hconfig][7] [28]),
        .I5(\slvi[haddr] [28]),
        .O(\slvi[hsel][7]_INST_0_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][7]_INST_0_i_23 
       (.I0(\slvo[7][hconfig][7] [8]),
        .I1(\slvo[7][hconfig][7] [24]),
        .I2(\slvi[haddr] [24]),
        .I3(\slvo[7][hconfig][7] [9]),
        .I4(\slvo[7][hconfig][7] [25]),
        .I5(\slvi[haddr] [25]),
        .O(\slvi[hsel][7]_INST_0_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D700D700D7D7D7)) 
    \slvi[hsel][7]_INST_0_i_24 
       (.I0(\slvo[7][hconfig][7] [5]),
        .I1(\slvo[7][hconfig][7] [21]),
        .I2(\slvi[haddr] [21]),
        .I3(\slvo[7][hconfig][7] [6]),
        .I4(\slvo[7][hconfig][7] [22]),
        .I5(\slvi[haddr] [22]),
        .O(\slvi[hsel][7]_INST_0_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000808030003000)) 
    \slvi[hsel][7]_INST_0_i_3 
       (.I0(hsel3),
        .I1(\slvo[7][hconfig][7] [0]),
        .I2(hsel2),
        .I3(hsel36_out),
        .I4(\slvi[hmbsel][2]_INST_0_i_9_n_0 ),
        .I5(\slvi[hmbsel][2]_INST_0_i_10_n_0 ),
        .O(\slvi[hsel][7]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][7]_INST_0_i_4 
       (.CI(slvi),
        .CO({hsel3,\slvi[hsel][7]_INST_0_i_4_n_1 ,\slvi[hsel][7]_INST_0_i_4_n_2 ,\slvi[hsel][7]_INST_0_i_4_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][7]_INST_0_i_7_n_0 ,\slvi[hsel][7]_INST_0_i_8_n_0 ,\slvi[hsel][7]_INST_0_i_9_n_0 ,\slvi[hsel][7]_INST_0_i_10_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \slvi[hsel][7]_INST_0_i_5 
       (.I0(\slvi[hsel][7]_INST_0_i_11_n_0 ),
        .I1(\slvi[hsel][7]_INST_0_i_12_n_0 ),
        .O(hsel2));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \slvi[hsel][7]_INST_0_i_6 
       (.CI(slvi),
        .CO({hsel36_out,\slvi[hsel][7]_INST_0_i_6_n_1 ,\slvi[hsel][7]_INST_0_i_6_n_2 ,\slvi[hsel][7]_INST_0_i_6_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({slvi,slvi,slvi,slvi}),
        .S({\slvi[hsel][7]_INST_0_i_13_n_0 ,\slvi[hsel][7]_INST_0_i_14_n_0 ,\slvi[hsel][7]_INST_0_i_15_n_0 ,\slvi[hsel][7]_INST_0_i_16_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][7]_INST_0_i_7 
       (.I0(\slvo[7][hconfig][7] [13]),
        .I1(\slvo[7][hconfig][7] [29]),
        .I2(\slvi[haddr] [17]),
        .I3(\slvi[hsel][7]_INST_0_i_17_n_0 ),
        .O(\slvi[hsel][7]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][7]_INST_0_i_8 
       (.I0(\slvo[7][hconfig][7] [10]),
        .I1(\slvo[7][hconfig][7] [26]),
        .I2(\slvi[haddr] [14]),
        .I3(\slvi[hsel][7]_INST_0_i_18_n_0 ),
        .O(\slvi[hsel][7]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hD700)) 
    \slvi[hsel][7]_INST_0_i_9 
       (.I0(\slvo[7][hconfig][7] [7]),
        .I1(\slvo[7][hconfig][7] [23]),
        .I2(\slvi[haddr] [11]),
        .I3(\slvi[hsel][7]_INST_0_i_19_n_0 ),
        .O(\slvi[hsel][7]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hsize][0]_INST_0 
       (.I0(\slvi[hsize][0]_INST_0_i_1_n_0 ),
        .I1(\slvi[hsize][0]_INST_0_i_2_n_0 ),
        .O(\slvi[hsize] [0]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hsize][0]_INST_0_i_1 
       (.I0(\msto[3][hsize] [0]),
        .I1(\msto[2][hsize] [0]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][hsize] [0]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][hsize] [0]),
        .O(\slvi[hsize][0]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hsize][0]_INST_0_i_2 
       (.I0(\msto[7][hsize] [0]),
        .I1(\msto[6][hsize] [0]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][hsize] [0]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][hsize] [0]),
        .O(\slvi[hsize][0]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hsize][1]_INST_0 
       (.I0(\slvi[hsize][1]_INST_0_i_1_n_0 ),
        .I1(\slvi[hsize][1]_INST_0_i_2_n_0 ),
        .O(\slvi[hsize] [1]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hsize][1]_INST_0_i_1 
       (.I0(\msto[3][hsize] [1]),
        .I1(\msto[2][hsize] [1]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][hsize] [1]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][hsize] [1]),
        .O(\slvi[hsize][1]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hsize][1]_INST_0_i_2 
       (.I0(\msto[7][hsize] [1]),
        .I1(\msto[6][hsize] [1]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][hsize] [1]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][hsize] [1]),
        .O(\slvi[hsize][1]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hsize][2]_INST_0 
       (.I0(\slvi[hsize][2]_INST_0_i_1_n_0 ),
        .I1(\slvi[hsize][2]_INST_0_i_2_n_0 ),
        .O(\slvi[hsize] [2]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hsize][2]_INST_0_i_1 
       (.I0(\msto[3][hsize] [2]),
        .I1(\msto[2][hsize] [2]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][hsize] [2]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][hsize] [2]),
        .O(\slvi[hsize][2]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hsize][2]_INST_0_i_2 
       (.I0(\msto[7][hsize] [2]),
        .I1(\msto[6][hsize] [2]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][hsize] [2]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][hsize] [2]),
        .O(\slvi[hsize][2]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[htrans][0]_INST_0 
       (.I0(\slvi[htrans][0]_INST_0_i_1_n_0 ),
        .I1(\slvi[htrans][0]_INST_0_i_2_n_0 ),
        .O(\slvi[htrans] [0]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[htrans][0]_INST_0_i_1 
       (.I0(\msto[3][htrans] [0]),
        .I1(\msto[2][htrans] [0]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][htrans] [0]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][htrans] [0]),
        .O(\slvi[htrans][0]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[htrans][0]_INST_0_i_2 
       (.I0(\msto[7][htrans] [0]),
        .I1(\msto[6][htrans] [0]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][htrans] [0]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][htrans] [0]),
        .O(\slvi[htrans][0]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[htrans][1]_INST_0 
       (.I0(\slvi[htrans][1]_INST_0_i_1_n_0 ),
        .I1(\slvi[htrans][1]_INST_0_i_2_n_0 ),
        .O(\slvi[htrans] [1]),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[htrans][1]_INST_0_i_1 
       (.I0(\msto[3][htrans] [1]),
        .I1(\msto[2][htrans] [1]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][htrans] [1]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][htrans] [1]),
        .O(\slvi[htrans][1]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[htrans][1]_INST_0_i_2 
       (.I0(\msto[7][htrans] [1]),
        .I1(\msto[6][htrans] [1]),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][htrans] [1]),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][htrans] [1]),
        .O(\slvi[htrans][1]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][0]_INST_0 
       (.I0(\slvi[hwdata][0]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][0]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [0]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][0]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [0]),
        .I1(\msto[2][hwdata] [0]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [0]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [0]),
        .O(\slvi[hwdata][0]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][0]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [0]),
        .I1(\msto[6][hwdata] [0]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [0]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [0]),
        .O(\slvi[hwdata][0]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][10]_INST_0 
       (.I0(\slvi[hwdata][10]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][10]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [10]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][10]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [10]),
        .I1(\msto[2][hwdata] [10]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [10]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [10]),
        .O(\slvi[hwdata][10]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][10]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [10]),
        .I1(\msto[6][hwdata] [10]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [10]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [10]),
        .O(\slvi[hwdata][10]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][11]_INST_0 
       (.I0(\slvi[hwdata][11]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][11]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [11]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][11]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [11]),
        .I1(\msto[2][hwdata] [11]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [11]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [11]),
        .O(\slvi[hwdata][11]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][11]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [11]),
        .I1(\msto[6][hwdata] [11]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [11]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [11]),
        .O(\slvi[hwdata][11]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][12]_INST_0 
       (.I0(\slvi[hwdata][12]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][12]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [12]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][12]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [12]),
        .I1(\msto[2][hwdata] [12]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [12]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [12]),
        .O(\slvi[hwdata][12]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][12]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [12]),
        .I1(\msto[6][hwdata] [12]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [12]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [12]),
        .O(\slvi[hwdata][12]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][13]_INST_0 
       (.I0(\slvi[hwdata][13]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][13]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [13]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][13]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [13]),
        .I1(\msto[2][hwdata] [13]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [13]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [13]),
        .O(\slvi[hwdata][13]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][13]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [13]),
        .I1(\msto[6][hwdata] [13]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [13]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [13]),
        .O(\slvi[hwdata][13]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][14]_INST_0 
       (.I0(\slvi[hwdata][14]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][14]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [14]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][14]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [14]),
        .I1(\msto[2][hwdata] [14]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [14]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [14]),
        .O(\slvi[hwdata][14]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][14]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [14]),
        .I1(\msto[6][hwdata] [14]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [14]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [14]),
        .O(\slvi[hwdata][14]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][15]_INST_0 
       (.I0(\slvi[hwdata][15]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][15]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [15]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][15]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [15]),
        .I1(\msto[2][hwdata] [15]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [15]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [15]),
        .O(\slvi[hwdata][15]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][15]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [15]),
        .I1(\msto[6][hwdata] [15]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [15]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [15]),
        .O(\slvi[hwdata][15]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][16]_INST_0 
       (.I0(\slvi[hwdata][16]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][16]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [16]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][16]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [16]),
        .I1(\msto[2][hwdata] [16]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [16]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [16]),
        .O(\slvi[hwdata][16]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][16]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [16]),
        .I1(\msto[6][hwdata] [16]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [16]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [16]),
        .O(\slvi[hwdata][16]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][17]_INST_0 
       (.I0(\slvi[hwdata][17]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][17]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [17]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][17]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [17]),
        .I1(\msto[2][hwdata] [17]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [17]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [17]),
        .O(\slvi[hwdata][17]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][17]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [17]),
        .I1(\msto[6][hwdata] [17]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [17]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [17]),
        .O(\slvi[hwdata][17]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][18]_INST_0 
       (.I0(\slvi[hwdata][18]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][18]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [18]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][18]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [18]),
        .I1(\msto[2][hwdata] [18]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [18]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [18]),
        .O(\slvi[hwdata][18]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][18]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [18]),
        .I1(\msto[6][hwdata] [18]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [18]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [18]),
        .O(\slvi[hwdata][18]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][19]_INST_0 
       (.I0(\slvi[hwdata][19]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][19]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [19]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][19]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [19]),
        .I1(\msto[2][hwdata] [19]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [19]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [19]),
        .O(\slvi[hwdata][19]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][19]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [19]),
        .I1(\msto[6][hwdata] [19]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [19]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [19]),
        .O(\slvi[hwdata][19]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][1]_INST_0 
       (.I0(\slvi[hwdata][1]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][1]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [1]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][1]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [1]),
        .I1(\msto[2][hwdata] [1]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [1]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [1]),
        .O(\slvi[hwdata][1]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][1]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [1]),
        .I1(\msto[6][hwdata] [1]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [1]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [1]),
        .O(\slvi[hwdata][1]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][20]_INST_0 
       (.I0(\slvi[hwdata][20]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][20]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [20]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][20]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [20]),
        .I1(\msto[2][hwdata] [20]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [20]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [20]),
        .O(\slvi[hwdata][20]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][20]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [20]),
        .I1(\msto[6][hwdata] [20]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [20]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [20]),
        .O(\slvi[hwdata][20]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][21]_INST_0 
       (.I0(\slvi[hwdata][21]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][21]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [21]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][21]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [21]),
        .I1(\msto[2][hwdata] [21]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [21]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [21]),
        .O(\slvi[hwdata][21]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][21]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [21]),
        .I1(\msto[6][hwdata] [21]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [21]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [21]),
        .O(\slvi[hwdata][21]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][22]_INST_0 
       (.I0(\slvi[hwdata][22]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][22]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [22]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][22]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [22]),
        .I1(\msto[2][hwdata] [22]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [22]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [22]),
        .O(\slvi[hwdata][22]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][22]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [22]),
        .I1(\msto[6][hwdata] [22]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [22]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [22]),
        .O(\slvi[hwdata][22]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][23]_INST_0 
       (.I0(\slvi[hwdata][23]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][23]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [23]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][23]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [23]),
        .I1(\msto[2][hwdata] [23]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [23]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [23]),
        .O(\slvi[hwdata][23]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][23]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [23]),
        .I1(\msto[6][hwdata] [23]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [23]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [23]),
        .O(\slvi[hwdata][23]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][24]_INST_0 
       (.I0(\slvi[hwdata][24]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][24]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [24]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][24]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [24]),
        .I1(\msto[2][hwdata] [24]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [24]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [24]),
        .O(\slvi[hwdata][24]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][24]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [24]),
        .I1(\msto[6][hwdata] [24]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [24]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [24]),
        .O(\slvi[hwdata][24]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][25]_INST_0 
       (.I0(\slvi[hwdata][25]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][25]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [25]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][25]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [25]),
        .I1(\msto[2][hwdata] [25]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [25]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [25]),
        .O(\slvi[hwdata][25]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][25]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [25]),
        .I1(\msto[6][hwdata] [25]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [25]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [25]),
        .O(\slvi[hwdata][25]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][26]_INST_0 
       (.I0(\slvi[hwdata][26]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][26]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [26]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][26]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [26]),
        .I1(\msto[2][hwdata] [26]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [26]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [26]),
        .O(\slvi[hwdata][26]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][26]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [26]),
        .I1(\msto[6][hwdata] [26]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [26]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [26]),
        .O(\slvi[hwdata][26]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][27]_INST_0 
       (.I0(\slvi[hwdata][27]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][27]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [27]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][27]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [27]),
        .I1(\msto[2][hwdata] [27]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [27]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [27]),
        .O(\slvi[hwdata][27]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][27]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [27]),
        .I1(\msto[6][hwdata] [27]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [27]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [27]),
        .O(\slvi[hwdata][27]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][28]_INST_0 
       (.I0(\slvi[hwdata][28]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][28]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [28]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][28]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [28]),
        .I1(\msto[2][hwdata] [28]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [28]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [28]),
        .O(\slvi[hwdata][28]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][28]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [28]),
        .I1(\msto[6][hwdata] [28]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [28]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [28]),
        .O(\slvi[hwdata][28]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][29]_INST_0 
       (.I0(\slvi[hwdata][29]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][29]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [29]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][29]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [29]),
        .I1(\msto[2][hwdata] [29]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [29]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [29]),
        .O(\slvi[hwdata][29]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][29]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [29]),
        .I1(\msto[6][hwdata] [29]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [29]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [29]),
        .O(\slvi[hwdata][29]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][2]_INST_0 
       (.I0(\slvi[hwdata][2]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][2]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [2]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][2]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [2]),
        .I1(\msto[2][hwdata] [2]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [2]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [2]),
        .O(\slvi[hwdata][2]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][2]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [2]),
        .I1(\msto[6][hwdata] [2]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [2]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [2]),
        .O(\slvi[hwdata][2]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][30]_INST_0 
       (.I0(\slvi[hwdata][30]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][30]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [30]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][30]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [30]),
        .I1(\msto[2][hwdata] [30]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [30]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [30]),
        .O(\slvi[hwdata][30]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][30]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [30]),
        .I1(\msto[6][hwdata] [30]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [30]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [30]),
        .O(\slvi[hwdata][30]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][31]_INST_0 
       (.I0(\slvi[hwdata][31]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][31]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [31]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][31]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [31]),
        .I1(\msto[2][hwdata] [31]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [31]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [31]),
        .O(\slvi[hwdata][31]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][31]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [31]),
        .I1(\msto[6][hwdata] [31]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [31]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [31]),
        .O(\slvi[hwdata][31]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][3]_INST_0 
       (.I0(\slvi[hwdata][3]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][3]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [3]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][3]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [3]),
        .I1(\msto[2][hwdata] [3]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [3]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [3]),
        .O(\slvi[hwdata][3]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][3]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [3]),
        .I1(\msto[6][hwdata] [3]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [3]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [3]),
        .O(\slvi[hwdata][3]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][4]_INST_0 
       (.I0(\slvi[hwdata][4]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][4]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [4]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][4]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [4]),
        .I1(\msto[2][hwdata] [4]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [4]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [4]),
        .O(\slvi[hwdata][4]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][4]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [4]),
        .I1(\msto[6][hwdata] [4]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [4]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [4]),
        .O(\slvi[hwdata][4]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][5]_INST_0 
       (.I0(\slvi[hwdata][5]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][5]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [5]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][5]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [5]),
        .I1(\msto[2][hwdata] [5]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [5]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [5]),
        .O(\slvi[hwdata][5]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][5]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [5]),
        .I1(\msto[6][hwdata] [5]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [5]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [5]),
        .O(\slvi[hwdata][5]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][6]_INST_0 
       (.I0(\slvi[hwdata][6]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][6]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [6]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][6]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [6]),
        .I1(\msto[2][hwdata] [6]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [6]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [6]),
        .O(\slvi[hwdata][6]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][6]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [6]),
        .I1(\msto[6][hwdata] [6]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [6]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [6]),
        .O(\slvi[hwdata][6]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][7]_INST_0 
       (.I0(\slvi[hwdata][7]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][7]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [7]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][7]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [7]),
        .I1(\msto[2][hwdata] [7]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [7]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [7]),
        .O(\slvi[hwdata][7]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][7]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [7]),
        .I1(\msto[6][hwdata] [7]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [7]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [7]),
        .O(\slvi[hwdata][7]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][8]_INST_0 
       (.I0(\slvi[hwdata][8]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][8]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [8]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][8]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [8]),
        .I1(\msto[2][hwdata] [8]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [8]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [8]),
        .O(\slvi[hwdata][8]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][8]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [8]),
        .I1(\msto[6][hwdata] [8]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [8]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [8]),
        .O(\slvi[hwdata][8]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwdata][9]_INST_0 
       (.I0(\slvi[hwdata][9]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwdata][9]_INST_0_i_2_n_0 ),
        .O(\slvi[hwdata] [9]),
        .S(\syncrregs.r_reg[hmasterd]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][9]_INST_0_i_1 
       (.I0(\msto[3][hwdata] [9]),
        .I1(\msto[2][hwdata] [9]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[1][hwdata] [9]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[0][hwdata] [9]),
        .O(\slvi[hwdata][9]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwdata][9]_INST_0_i_2 
       (.I0(\msto[7][hwdata] [9]),
        .I1(\msto[6][hwdata] [9]),
        .I2(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I3(\msto[5][hwdata] [9]),
        .I4(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I5(\msto[4][hwdata] [9]),
        .O(\slvi[hwdata][9]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \slvi[hwrite]_INST_0 
       (.I0(\slvi[hwrite]_INST_0_i_1_n_0 ),
        .I1(\slvi[hwrite]_INST_0_i_2_n_0 ),
        .O(\slvi[hwrite] ),
        .S(\^slvi[hmaster] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwrite]_INST_0_i_1 
       (.I0(\msto[3][hwrite] ),
        .I1(\msto[2][hwrite] ),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[1][hwrite] ),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[0][hwrite] ),
        .O(\slvi[hwrite]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \slvi[hwrite]_INST_0_i_2 
       (.I0(\msto[7][hwrite] ),
        .I1(\msto[6][hwrite] ),
        .I2(\^slvi[hmaster] [1]),
        .I3(\msto[5][hwrite] ),
        .I4(\^slvi[hmaster] [0]),
        .I5(\msto[4][hwrite] ),
        .O(\slvi[hwrite]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \slvi[testin][2]_INST_0 
       (.I0(testen),
        .I1(scanen),
        .O(\^slvi[testin] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \syncrregs.r[defslv]_i_1 
       (.I0(p_14_out),
        .I1(\^slvi[hsel] [0]),
        .I2(hsel1192_out),
        .I3(p_6_out),
        .I4(p_11_out),
        .O(p_185_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \syncrregs.r[hmaster][0]_i_1 
       (.I0(\syncrregs.r[hmaster][0]_i_2_n_0 ),
        .I1(rst),
        .O(\syncrregs.r ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAACAAAAAAAAAAAAA)) 
    \syncrregs.r[hmaster][0]_i_2 
       (.I0(\^slvi[hmaster] [0]),
        .I1(\msti[hgrant][0]_INST_0_i_10_n_0 ),
        .I2(\msti[hgrant][0]_INST_0_i_6_n_0 ),
        .I3(\msti[hgrant][0]_INST_0_i_8_n_0 ),
        .I4(\slvi[hready] ),
        .I5(arb1_out),
        .O(\syncrregs.r[hmaster][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \syncrregs.r[hmaster][1]_i_1 
       (.I0(\syncrregs.r[hmaster][1]_i_2_n_0 ),
        .I1(rst),
        .O(\syncrregs.r[hmaster][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAACAAAAAAAAAAAAA)) 
    \syncrregs.r[hmaster][1]_i_2 
       (.I0(\^slvi[hmaster] [1]),
        .I1(\msti[hgrant][0]_INST_0_i_5_n_0 ),
        .I2(\msti[hgrant][0]_INST_0_i_6_n_0 ),
        .I3(\msti[hgrant][0]_INST_0_i_8_n_0 ),
        .I4(\slvi[hready] ),
        .I5(arb1_out),
        .O(\syncrregs.r[hmaster][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \syncrregs.r[hmaster][2]_i_1 
       (.I0(\syncrregs.r[hmaster][2]_i_2_n_0 ),
        .I1(rst),
        .O(\syncrregs.r[hmaster][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAACAAAAAAAAAAAAA)) 
    \syncrregs.r[hmaster][2]_i_2 
       (.I0(\^slvi[hmaster] [2]),
        .I1(\msti[hgrant][0]_INST_0_i_12_n_0 ),
        .I2(\msti[hgrant][0]_INST_0_i_6_n_0 ),
        .I3(\msti[hgrant][0]_INST_0_i_8_n_0 ),
        .I4(\slvi[hready] ),
        .I5(arb1_out),
        .O(\syncrregs.r[hmaster][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000F400)) 
    \syncrregs.r[hmasterlock]_i_1 
       (.I0(\slvi[hready] ),
        .I1(\slvi[hmastlock] ),
        .I2(\syncrregs.r_reg[hmasterlock]_i_2_n_0 ),
        .I3(rst),
        .I4(v),
        .O(\syncrregs.r[hmasterlock]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000090000000)) 
    \syncrregs.r[hmasterlock]_i_3 
       (.I0(\syncrregs.r[hmaster][0]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hmasterd]__0 [0]),
        .I2(\syncrregs.r[hmasterlock]_i_6_n_0 ),
        .I3(\syncrregs.r[hmasterlock]_i_7_n_0 ),
        .I4(p_0_in186_in),
        .I5(\syncrregs.r_reg[hmasterlockd]__0 ),
        .O(v));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hmasterlock]_i_4 
       (.I0(\msto[3][hlock] ),
        .I1(\msto[2][hlock] ),
        .I2(\syncrregs.r[hmaster][1]_i_2_n_0 ),
        .I3(\msto[1][hlock] ),
        .I4(\syncrregs.r[hmaster][0]_i_2_n_0 ),
        .I5(\msto[0][hlock] ),
        .O(\syncrregs.r[hmasterlock]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hmasterlock]_i_5 
       (.I0(\msto[7][hlock] ),
        .I1(\msto[6][hlock] ),
        .I2(\syncrregs.r[hmaster][1]_i_2_n_0 ),
        .I3(\msto[5][hlock] ),
        .I4(\syncrregs.r[hmaster][0]_i_2_n_0 ),
        .I5(\msto[4][hlock] ),
        .O(\syncrregs.r[hmasterlock]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAA9AA56555555)) 
    \syncrregs.r[hmasterlock]_i_6 
       (.I0(\syncrregs.r_reg[hmasterd]__0 [2]),
        .I1(\syncrregs.r[hmasterlock]_i_8_n_0 ),
        .I2(\msti[hgrant][0]_INST_0_i_8_n_0 ),
        .I3(\msti[hgrant][0]_INST_0_i_6_n_0 ),
        .I4(\msti[hgrant][0]_INST_0_i_12_n_0 ),
        .I5(\^slvi[hmaster] [2]),
        .O(\syncrregs.r[hmasterlock]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAA9AA56555555)) 
    \syncrregs.r[hmasterlock]_i_7 
       (.I0(\syncrregs.r_reg[hmasterd]__0 [1]),
        .I1(\syncrregs.r[hmasterlock]_i_8_n_0 ),
        .I2(\msti[hgrant][0]_INST_0_i_8_n_0 ),
        .I3(\msti[hgrant][0]_INST_0_i_6_n_0 ),
        .I4(\msti[hgrant][0]_INST_0_i_5_n_0 ),
        .I5(\^slvi[hmaster] [1]),
        .O(\syncrregs.r[hmasterlock]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \syncrregs.r[hmasterlock]_i_8 
       (.I0(\slvi[hready] ),
        .I1(arb1_out),
        .O(\syncrregs.r[hmasterlock]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0B08)) 
    \syncrregs.r[hmasterlockd]_i_1 
       (.I0(\slvi[hmastlock] ),
        .I1(\slvi[hready] ),
        .I2(v),
        .I3(\syncrregs.r_reg[hmasterlockd]__0 ),
        .O(\syncrregs.r[hmasterlockd]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][0]_i_2 
       (.I0(\msto[3][hconfig][0] [0]),
        .I1(\msto[2][hconfig][0] [0]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [0]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [0]),
        .O(\syncrregs.r[hrdatam][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][0]_i_3 
       (.I0(\msto[7][hconfig][0] [0]),
        .I1(\msto[6][hconfig][0] [0]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [0]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [0]),
        .O(\syncrregs.r[hrdatam][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][10]_i_2 
       (.I0(\msto[3][hconfig][0] [10]),
        .I1(\msto[2][hconfig][0] [10]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [10]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [10]),
        .O(\syncrregs.r[hrdatam][10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][10]_i_3 
       (.I0(\msto[7][hconfig][0] [10]),
        .I1(\msto[6][hconfig][0] [10]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [10]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [10]),
        .O(\syncrregs.r[hrdatam][10]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][11]_i_2 
       (.I0(\msto[3][hconfig][0] [11]),
        .I1(\msto[2][hconfig][0] [11]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [11]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [11]),
        .O(\syncrregs.r[hrdatam][11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][11]_i_3 
       (.I0(\msto[7][hconfig][0] [11]),
        .I1(\msto[6][hconfig][0] [11]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [11]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [11]),
        .O(\syncrregs.r[hrdatam][11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][12]_i_2 
       (.I0(\msto[3][hconfig][0] [12]),
        .I1(\msto[2][hconfig][0] [12]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [12]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [12]),
        .O(\syncrregs.r[hrdatam][12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][12]_i_3 
       (.I0(\msto[7][hconfig][0] [12]),
        .I1(\msto[6][hconfig][0] [12]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [12]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [12]),
        .O(\syncrregs.r[hrdatam][12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][13]_i_2 
       (.I0(\msto[3][hconfig][0] [13]),
        .I1(\msto[2][hconfig][0] [13]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [13]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [13]),
        .O(\syncrregs.r[hrdatam][13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][13]_i_3 
       (.I0(\msto[7][hconfig][0] [13]),
        .I1(\msto[6][hconfig][0] [13]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [13]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [13]),
        .O(\syncrregs.r[hrdatam][13]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][14]_i_2 
       (.I0(\msto[3][hconfig][0] [14]),
        .I1(\msto[2][hconfig][0] [14]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [14]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [14]),
        .O(\syncrregs.r[hrdatam][14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][14]_i_3 
       (.I0(\msto[7][hconfig][0] [14]),
        .I1(\msto[6][hconfig][0] [14]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [14]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [14]),
        .O(\syncrregs.r[hrdatam][14]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][15]_i_2 
       (.I0(\msto[3][hconfig][0] [15]),
        .I1(\msto[2][hconfig][0] [15]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [15]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [15]),
        .O(\syncrregs.r[hrdatam][15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][15]_i_3 
       (.I0(\msto[7][hconfig][0] [15]),
        .I1(\msto[6][hconfig][0] [15]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [15]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [15]),
        .O(\syncrregs.r[hrdatam][15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][16]_i_2 
       (.I0(\msto[3][hconfig][0] [16]),
        .I1(\msto[2][hconfig][0] [16]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [16]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [16]),
        .O(\syncrregs.r[hrdatam][16]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][16]_i_3 
       (.I0(\msto[7][hconfig][0] [16]),
        .I1(\msto[6][hconfig][0] [16]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [16]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [16]),
        .O(\syncrregs.r[hrdatam][16]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][17]_i_2 
       (.I0(\msto[3][hconfig][0] [17]),
        .I1(\msto[2][hconfig][0] [17]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [17]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [17]),
        .O(\syncrregs.r[hrdatam][17]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][17]_i_3 
       (.I0(\msto[7][hconfig][0] [17]),
        .I1(\msto[6][hconfig][0] [17]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [17]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [17]),
        .O(\syncrregs.r[hrdatam][17]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][18]_i_2 
       (.I0(\msto[3][hconfig][0] [18]),
        .I1(\msto[2][hconfig][0] [18]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [18]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [18]),
        .O(\syncrregs.r[hrdatam][18]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][18]_i_3 
       (.I0(\msto[7][hconfig][0] [18]),
        .I1(\msto[6][hconfig][0] [18]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [18]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [18]),
        .O(\syncrregs.r[hrdatam][18]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][19]_i_2 
       (.I0(\msto[3][hconfig][0] [19]),
        .I1(\msto[2][hconfig][0] [19]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [19]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [19]),
        .O(\syncrregs.r[hrdatam][19]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][19]_i_3 
       (.I0(\msto[7][hconfig][0] [19]),
        .I1(\msto[6][hconfig][0] [19]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [19]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [19]),
        .O(\syncrregs.r[hrdatam][19]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][1]_i_2 
       (.I0(\msto[3][hconfig][0] [1]),
        .I1(\msto[2][hconfig][0] [1]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [1]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [1]),
        .O(\syncrregs.r[hrdatam][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][1]_i_3 
       (.I0(\msto[7][hconfig][0] [1]),
        .I1(\msto[6][hconfig][0] [1]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [1]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [1]),
        .O(\syncrregs.r[hrdatam][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][20]_i_2 
       (.I0(\msto[3][hconfig][0] [20]),
        .I1(\msto[2][hconfig][0] [20]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [20]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [20]),
        .O(\syncrregs.r[hrdatam][20]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][20]_i_3 
       (.I0(\msto[7][hconfig][0] [20]),
        .I1(\msto[6][hconfig][0] [20]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [20]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [20]),
        .O(\syncrregs.r[hrdatam][20]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][21]_i_2 
       (.I0(\msto[3][hconfig][0] [21]),
        .I1(\msto[2][hconfig][0] [21]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [21]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [21]),
        .O(\syncrregs.r[hrdatam][21]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][21]_i_3 
       (.I0(\msto[7][hconfig][0] [21]),
        .I1(\msto[6][hconfig][0] [21]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [21]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [21]),
        .O(\syncrregs.r[hrdatam][21]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][22]_i_2 
       (.I0(\msto[3][hconfig][0] [22]),
        .I1(\msto[2][hconfig][0] [22]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [22]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [22]),
        .O(\syncrregs.r[hrdatam][22]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][22]_i_3 
       (.I0(\msto[7][hconfig][0] [22]),
        .I1(\msto[6][hconfig][0] [22]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [22]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [22]),
        .O(\syncrregs.r[hrdatam][22]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][23]_i_2 
       (.I0(\msto[3][hconfig][0] [23]),
        .I1(\msto[2][hconfig][0] [23]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [23]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [23]),
        .O(\syncrregs.r[hrdatam][23]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][23]_i_3 
       (.I0(\msto[7][hconfig][0] [23]),
        .I1(\msto[6][hconfig][0] [23]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [23]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [23]),
        .O(\syncrregs.r[hrdatam][23]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][24]_i_2 
       (.I0(\msto[3][hconfig][0] [24]),
        .I1(\msto[2][hconfig][0] [24]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [24]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [24]),
        .O(\syncrregs.r[hrdatam][24]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][24]_i_3 
       (.I0(\msto[7][hconfig][0] [24]),
        .I1(\msto[6][hconfig][0] [24]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [24]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [24]),
        .O(\syncrregs.r[hrdatam][24]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][25]_i_2 
       (.I0(\msto[3][hconfig][0] [25]),
        .I1(\msto[2][hconfig][0] [25]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [25]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [25]),
        .O(\syncrregs.r[hrdatam][25]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][25]_i_3 
       (.I0(\msto[7][hconfig][0] [25]),
        .I1(\msto[6][hconfig][0] [25]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [25]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [25]),
        .O(\syncrregs.r[hrdatam][25]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][26]_i_2 
       (.I0(\msto[3][hconfig][0] [26]),
        .I1(\msto[2][hconfig][0] [26]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [26]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [26]),
        .O(\syncrregs.r[hrdatam][26]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][26]_i_3 
       (.I0(\msto[7][hconfig][0] [26]),
        .I1(\msto[6][hconfig][0] [26]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [26]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [26]),
        .O(\syncrregs.r[hrdatam][26]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][27]_i_2 
       (.I0(\msto[3][hconfig][0] [27]),
        .I1(\msto[2][hconfig][0] [27]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [27]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [27]),
        .O(\syncrregs.r[hrdatam][27]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][27]_i_3 
       (.I0(\msto[7][hconfig][0] [27]),
        .I1(\msto[6][hconfig][0] [27]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [27]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [27]),
        .O(\syncrregs.r[hrdatam][27]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][28]_i_2 
       (.I0(\msto[3][hconfig][0] [28]),
        .I1(\msto[2][hconfig][0] [28]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [28]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [28]),
        .O(\syncrregs.r[hrdatam][28]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][28]_i_3 
       (.I0(\msto[7][hconfig][0] [28]),
        .I1(\msto[6][hconfig][0] [28]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [28]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [28]),
        .O(\syncrregs.r[hrdatam][28]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][29]_i_2 
       (.I0(\msto[3][hconfig][0] [29]),
        .I1(\msto[2][hconfig][0] [29]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [29]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [29]),
        .O(\syncrregs.r[hrdatam][29]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][29]_i_3 
       (.I0(\msto[7][hconfig][0] [29]),
        .I1(\msto[6][hconfig][0] [29]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [29]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [29]),
        .O(\syncrregs.r[hrdatam][29]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][2]_i_2 
       (.I0(\msto[3][hconfig][0] [2]),
        .I1(\msto[2][hconfig][0] [2]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [2]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [2]),
        .O(\syncrregs.r[hrdatam][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][2]_i_3 
       (.I0(\msto[7][hconfig][0] [2]),
        .I1(\msto[6][hconfig][0] [2]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [2]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [2]),
        .O(\syncrregs.r[hrdatam][2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][30]_i_2 
       (.I0(\msto[3][hconfig][0] [30]),
        .I1(\msto[2][hconfig][0] [30]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [30]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [30]),
        .O(\syncrregs.r[hrdatam][30]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][30]_i_3 
       (.I0(\msto[7][hconfig][0] [30]),
        .I1(\msto[6][hconfig][0] [30]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [30]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [30]),
        .O(\syncrregs.r[hrdatam][30]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \syncrregs.r[hrdatam][31]_i_1 
       (.I0(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I1(\syncrregs.r_reg[haddr_n_0_][2] ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(sel0[5]),
        .I4(sel0[4]),
        .I5(sel0[6]),
        .O(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][31]_i_3 
       (.I0(\msto[3][hconfig][0] [31]),
        .I1(\msto[2][hconfig][0] [31]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [31]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [31]),
        .O(\syncrregs.r[hrdatam][31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][31]_i_4 
       (.I0(\msto[7][hconfig][0] [31]),
        .I1(\msto[6][hconfig][0] [31]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [31]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [31]),
        .O(\syncrregs.r[hrdatam][31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][3]_i_2 
       (.I0(\msto[3][hconfig][0] [3]),
        .I1(\msto[2][hconfig][0] [3]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [3]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [3]),
        .O(\syncrregs.r[hrdatam][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][3]_i_3 
       (.I0(\msto[7][hconfig][0] [3]),
        .I1(\msto[6][hconfig][0] [3]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [3]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [3]),
        .O(\syncrregs.r[hrdatam][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][4]_i_2 
       (.I0(\msto[3][hconfig][0] [4]),
        .I1(\msto[2][hconfig][0] [4]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [4]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [4]),
        .O(\syncrregs.r[hrdatam][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][4]_i_3 
       (.I0(\msto[7][hconfig][0] [4]),
        .I1(\msto[6][hconfig][0] [4]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [4]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [4]),
        .O(\syncrregs.r[hrdatam][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][5]_i_2 
       (.I0(\msto[3][hconfig][0] [5]),
        .I1(\msto[2][hconfig][0] [5]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [5]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [5]),
        .O(\syncrregs.r[hrdatam][5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][5]_i_3 
       (.I0(\msto[7][hconfig][0] [5]),
        .I1(\msto[6][hconfig][0] [5]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [5]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [5]),
        .O(\syncrregs.r[hrdatam][5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][6]_i_2 
       (.I0(\msto[3][hconfig][0] [6]),
        .I1(\msto[2][hconfig][0] [6]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [6]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [6]),
        .O(\syncrregs.r[hrdatam][6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][6]_i_3 
       (.I0(\msto[7][hconfig][0] [6]),
        .I1(\msto[6][hconfig][0] [6]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [6]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [6]),
        .O(\syncrregs.r[hrdatam][6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][7]_i_2 
       (.I0(\msto[3][hconfig][0] [7]),
        .I1(\msto[2][hconfig][0] [7]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [7]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [7]),
        .O(\syncrregs.r[hrdatam][7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][7]_i_3 
       (.I0(\msto[7][hconfig][0] [7]),
        .I1(\msto[6][hconfig][0] [7]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [7]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [7]),
        .O(\syncrregs.r[hrdatam][7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][8]_i_2 
       (.I0(\msto[3][hconfig][0] [8]),
        .I1(\msto[2][hconfig][0] [8]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [8]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [8]),
        .O(\syncrregs.r[hrdatam][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][8]_i_3 
       (.I0(\msto[7][hconfig][0] [8]),
        .I1(\msto[6][hconfig][0] [8]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [8]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [8]),
        .O(\syncrregs.r[hrdatam][8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][9]_i_2 
       (.I0(\msto[3][hconfig][0] [9]),
        .I1(\msto[2][hconfig][0] [9]),
        .I2(sel0[2]),
        .I3(\msto[1][hconfig][0] [9]),
        .I4(sel0[1]),
        .I5(\msto[0][hconfig][0] [9]),
        .O(\syncrregs.r[hrdatam][9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatam][9]_i_3 
       (.I0(\msto[7][hconfig][0] [9]),
        .I1(\msto[6][hconfig][0] [9]),
        .I2(sel0[2]),
        .I3(\msto[5][hconfig][0] [9]),
        .I4(sel0[1]),
        .I5(\msto[4][hconfig][0] [9]),
        .O(\syncrregs.r[hrdatam][9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][0]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][0]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][0]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][0]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][0]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][0]_i_14 
       (.I0(\slvo[3][hconfig][6] [0]),
        .I1(\slvo[2][hconfig][6] [0]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][6] [0]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][6] [0]),
        .O(\syncrregs.r[hrdatas][0]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][0]_i_15 
       (.I0(\slvo[7][hconfig][6] [0]),
        .I1(\slvo[6][hconfig][6] [0]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][6] [0]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][6] [0]),
        .O(\syncrregs.r[hrdatas][0]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][0]_i_16 
       (.I0(\slvo[3][hconfig][7] [0]),
        .I1(\slvo[2][hconfig][7] [0]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][7] [0]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][7] [0]),
        .O(\syncrregs.r[hrdatas][0]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][0]_i_17 
       (.I0(\slvo[7][hconfig][7] [0]),
        .I1(\slvo[6][hconfig][7] [0]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][7] [0]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][7] [0]),
        .O(\syncrregs.r[hrdatas][0]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][0]_i_18 
       (.I0(\slvo[3][hconfig][4] [0]),
        .I1(\slvo[2][hconfig][4] [0]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][4] [0]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][4] [0]),
        .O(\syncrregs.r[hrdatas][0]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][0]_i_19 
       (.I0(\slvo[7][hconfig][4] [0]),
        .I1(\slvo[6][hconfig][4] [0]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][4] [0]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][4] [0]),
        .O(\syncrregs.r[hrdatas][0]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][0]_i_20 
       (.I0(\slvo[3][hconfig][5] [0]),
        .I1(\slvo[2][hconfig][5] [0]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][5] [0]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][5] [0]),
        .O(\syncrregs.r[hrdatas][0]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][0]_i_21 
       (.I0(\slvo[7][hconfig][5] [0]),
        .I1(\slvo[6][hconfig][5] [0]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][5] [0]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][5] [0]),
        .O(\syncrregs.r[hrdatas][0]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][0]_i_22 
       (.I0(\slvo[3][hconfig][2] [0]),
        .I1(\slvo[2][hconfig][2] [0]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][2] [0]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][2] [0]),
        .O(\syncrregs.r[hrdatas][0]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][0]_i_23 
       (.I0(\slvo[7][hconfig][2] [0]),
        .I1(\slvo[6][hconfig][2] [0]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][2] [0]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][2] [0]),
        .O(\syncrregs.r[hrdatas][0]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][0]_i_24 
       (.I0(\slvo[3][hconfig][3] [0]),
        .I1(\slvo[2][hconfig][3] [0]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][3] [0]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][3] [0]),
        .O(\syncrregs.r[hrdatas][0]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][0]_i_25 
       (.I0(\slvo[7][hconfig][3] [0]),
        .I1(\slvo[6][hconfig][3] [0]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][3] [0]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][3] [0]),
        .O(\syncrregs.r[hrdatas][0]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][0]_i_26 
       (.I0(\slvo[3][hconfig][0] [0]),
        .I1(\slvo[2][hconfig][0] [0]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][0] [0]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][0] [0]),
        .O(\syncrregs.r[hrdatas][0]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][0]_i_27 
       (.I0(\slvo[7][hconfig][0] [0]),
        .I1(\slvo[6][hconfig][0] [0]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][0] [0]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][0] [0]),
        .O(\syncrregs.r[hrdatas][0]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][0]_i_28 
       (.I0(\slvo[3][hconfig][1] [0]),
        .I1(\slvo[2][hconfig][1] [0]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][1] [0]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][1] [0]),
        .O(\syncrregs.r[hrdatas][0]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][0]_i_29 
       (.I0(\slvo[7][hconfig][1] [0]),
        .I1(\slvo[6][hconfig][1] [0]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][1] [0]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][1] [0]),
        .O(\syncrregs.r[hrdatas][0]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][10]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][10]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][10]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][10]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][10]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][10]_i_14 
       (.I0(\slvo[3][hconfig][6] [10]),
        .I1(\slvo[2][hconfig][6] [10]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][6] [10]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][6] [10]),
        .O(\syncrregs.r[hrdatas][10]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][10]_i_15 
       (.I0(\slvo[7][hconfig][6] [10]),
        .I1(\slvo[6][hconfig][6] [10]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][6] [10]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][6] [10]),
        .O(\syncrregs.r[hrdatas][10]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][10]_i_16 
       (.I0(\slvo[3][hconfig][7] [10]),
        .I1(\slvo[2][hconfig][7] [10]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][7] [10]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][7] [10]),
        .O(\syncrregs.r[hrdatas][10]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][10]_i_17 
       (.I0(\slvo[7][hconfig][7] [10]),
        .I1(\slvo[6][hconfig][7] [10]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][7] [10]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][7] [10]),
        .O(\syncrregs.r[hrdatas][10]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][10]_i_18 
       (.I0(\slvo[3][hconfig][4] [10]),
        .I1(\slvo[2][hconfig][4] [10]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][4] [10]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][4] [10]),
        .O(\syncrregs.r[hrdatas][10]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][10]_i_19 
       (.I0(\slvo[7][hconfig][4] [10]),
        .I1(\slvo[6][hconfig][4] [10]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][4] [10]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][4] [10]),
        .O(\syncrregs.r[hrdatas][10]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][10]_i_20 
       (.I0(\slvo[3][hconfig][5] [10]),
        .I1(\slvo[2][hconfig][5] [10]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][5] [10]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][5] [10]),
        .O(\syncrregs.r[hrdatas][10]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][10]_i_21 
       (.I0(\slvo[7][hconfig][5] [10]),
        .I1(\slvo[6][hconfig][5] [10]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][5] [10]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][5] [10]),
        .O(\syncrregs.r[hrdatas][10]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][10]_i_22 
       (.I0(\slvo[3][hconfig][2] [10]),
        .I1(\slvo[2][hconfig][2] [10]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][2] [10]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][2] [10]),
        .O(\syncrregs.r[hrdatas][10]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][10]_i_23 
       (.I0(\slvo[7][hconfig][2] [10]),
        .I1(\slvo[6][hconfig][2] [10]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][2] [10]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][2] [10]),
        .O(\syncrregs.r[hrdatas][10]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][10]_i_24 
       (.I0(\slvo[3][hconfig][3] [10]),
        .I1(\slvo[2][hconfig][3] [10]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][3] [10]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][3] [10]),
        .O(\syncrregs.r[hrdatas][10]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][10]_i_25 
       (.I0(\slvo[7][hconfig][3] [10]),
        .I1(\slvo[6][hconfig][3] [10]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][3] [10]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][3] [10]),
        .O(\syncrregs.r[hrdatas][10]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][10]_i_26 
       (.I0(\slvo[3][hconfig][0] [10]),
        .I1(\slvo[2][hconfig][0] [10]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][0] [10]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][0] [10]),
        .O(\syncrregs.r[hrdatas][10]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][10]_i_27 
       (.I0(\slvo[7][hconfig][0] [10]),
        .I1(\slvo[6][hconfig][0] [10]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][0] [10]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][0] [10]),
        .O(\syncrregs.r[hrdatas][10]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][10]_i_28 
       (.I0(\slvo[3][hconfig][1] [10]),
        .I1(\slvo[2][hconfig][1] [10]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][1] [10]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][1] [10]),
        .O(\syncrregs.r[hrdatas][10]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][10]_i_29 
       (.I0(\slvo[7][hconfig][1] [10]),
        .I1(\slvo[6][hconfig][1] [10]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][1] [10]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][1] [10]),
        .O(\syncrregs.r[hrdatas][10]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][11]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][11]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][11]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][11]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][11]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][11]_i_14 
       (.I0(\slvo[3][hconfig][6] [11]),
        .I1(\slvo[2][hconfig][6] [11]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][6] [11]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][6] [11]),
        .O(\syncrregs.r[hrdatas][11]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][11]_i_15 
       (.I0(\slvo[7][hconfig][6] [11]),
        .I1(\slvo[6][hconfig][6] [11]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][6] [11]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][6] [11]),
        .O(\syncrregs.r[hrdatas][11]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][11]_i_16 
       (.I0(\slvo[3][hconfig][7] [11]),
        .I1(\slvo[2][hconfig][7] [11]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][7] [11]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][7] [11]),
        .O(\syncrregs.r[hrdatas][11]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][11]_i_17 
       (.I0(\slvo[7][hconfig][7] [11]),
        .I1(\slvo[6][hconfig][7] [11]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][7] [11]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][7] [11]),
        .O(\syncrregs.r[hrdatas][11]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][11]_i_18 
       (.I0(\slvo[3][hconfig][4] [11]),
        .I1(\slvo[2][hconfig][4] [11]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][4] [11]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][4] [11]),
        .O(\syncrregs.r[hrdatas][11]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][11]_i_19 
       (.I0(\slvo[7][hconfig][4] [11]),
        .I1(\slvo[6][hconfig][4] [11]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][4] [11]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][4] [11]),
        .O(\syncrregs.r[hrdatas][11]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][11]_i_20 
       (.I0(\slvo[3][hconfig][5] [11]),
        .I1(\slvo[2][hconfig][5] [11]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][5] [11]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][5] [11]),
        .O(\syncrregs.r[hrdatas][11]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][11]_i_21 
       (.I0(\slvo[7][hconfig][5] [11]),
        .I1(\slvo[6][hconfig][5] [11]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][5] [11]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][5] [11]),
        .O(\syncrregs.r[hrdatas][11]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][11]_i_22 
       (.I0(\slvo[3][hconfig][2] [11]),
        .I1(\slvo[2][hconfig][2] [11]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][2] [11]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][2] [11]),
        .O(\syncrregs.r[hrdatas][11]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][11]_i_23 
       (.I0(\slvo[7][hconfig][2] [11]),
        .I1(\slvo[6][hconfig][2] [11]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][2] [11]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][2] [11]),
        .O(\syncrregs.r[hrdatas][11]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][11]_i_24 
       (.I0(\slvo[3][hconfig][3] [11]),
        .I1(\slvo[2][hconfig][3] [11]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][3] [11]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][3] [11]),
        .O(\syncrregs.r[hrdatas][11]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][11]_i_25 
       (.I0(\slvo[7][hconfig][3] [11]),
        .I1(\slvo[6][hconfig][3] [11]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][3] [11]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][3] [11]),
        .O(\syncrregs.r[hrdatas][11]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][11]_i_26 
       (.I0(\slvo[3][hconfig][0] [11]),
        .I1(\slvo[2][hconfig][0] [11]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][0] [11]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][0] [11]),
        .O(\syncrregs.r[hrdatas][11]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][11]_i_27 
       (.I0(\slvo[7][hconfig][0] [11]),
        .I1(\slvo[6][hconfig][0] [11]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][0] [11]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][0] [11]),
        .O(\syncrregs.r[hrdatas][11]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][11]_i_28 
       (.I0(\slvo[3][hconfig][1] [11]),
        .I1(\slvo[2][hconfig][1] [11]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][1] [11]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][1] [11]),
        .O(\syncrregs.r[hrdatas][11]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][11]_i_29 
       (.I0(\slvo[7][hconfig][1] [11]),
        .I1(\slvo[6][hconfig][1] [11]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][1] [11]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][1] [11]),
        .O(\syncrregs.r[hrdatas][11]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \syncrregs.r[hrdatas][12]_i_1 
       (.I0(sel0[6]),
        .I1(\syncrregs.r[hrdatas][12]_i_3_n_0 ),
        .O(\v[hrdatas] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][12]_i_15 
       (.I0(\slvo[3][hconfig][3] [12]),
        .I1(\slvo[2][hconfig][3] [12]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][3] [12]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][3] [12]),
        .O(\syncrregs.r[hrdatas][12]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][12]_i_16 
       (.I0(\slvo[7][hconfig][3] [12]),
        .I1(\slvo[6][hconfig][3] [12]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][3] [12]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][3] [12]),
        .O(\syncrregs.r[hrdatas][12]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][12]_i_17 
       (.I0(\slvo[3][hconfig][2] [12]),
        .I1(\slvo[2][hconfig][2] [12]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][2] [12]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][2] [12]),
        .O(\syncrregs.r[hrdatas][12]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][12]_i_18 
       (.I0(\slvo[7][hconfig][2] [12]),
        .I1(\slvo[6][hconfig][2] [12]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][2] [12]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][2] [12]),
        .O(\syncrregs.r[hrdatas][12]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][12]_i_19 
       (.I0(\slvo[3][hconfig][1] [12]),
        .I1(\slvo[2][hconfig][1] [12]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][1] [12]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][1] [12]),
        .O(\syncrregs.r[hrdatas][12]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEE222E200000000)) 
    \syncrregs.r[hrdatas][12]_i_2 
       (.I0(\syncrregs.r[hrdatas][12]_i_4_n_0 ),
        .I1(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I2(\syncrregs.r_reg[hrdatas][12]_i_5_n_0 ),
        .I3(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I4(\syncrregs.r_reg[hrdatas][12]_i_6_n_0 ),
        .I5(p_179_out),
        .O(\syncrregs.r[hrdatas][12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][12]_i_20 
       (.I0(\slvo[7][hconfig][1] [12]),
        .I1(\slvo[6][hconfig][1] [12]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][1] [12]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][1] [12]),
        .O(\syncrregs.r[hrdatas][12]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][12]_i_21 
       (.I0(\slvo[3][hconfig][0] [12]),
        .I1(\slvo[2][hconfig][0] [12]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][0] [12]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][0] [12]),
        .O(\syncrregs.r[hrdatas][12]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][12]_i_22 
       (.I0(\slvo[7][hconfig][0] [12]),
        .I1(\slvo[6][hconfig][0] [12]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][0] [12]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][0] [12]),
        .O(\syncrregs.r[hrdatas][12]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][12]_i_23 
       (.I0(\slvo[3][hconfig][4] [12]),
        .I1(\slvo[2][hconfig][4] [12]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][4] [12]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][4] [12]),
        .O(\syncrregs.r[hrdatas][12]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][12]_i_24 
       (.I0(\slvo[7][hconfig][4] [12]),
        .I1(\slvo[6][hconfig][4] [12]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][4] [12]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][4] [12]),
        .O(\syncrregs.r[hrdatas][12]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][12]_i_25 
       (.I0(\slvo[3][hconfig][5] [12]),
        .I1(\slvo[2][hconfig][5] [12]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][5] [12]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][5] [12]),
        .O(\syncrregs.r[hrdatas][12]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][12]_i_26 
       (.I0(\slvo[7][hconfig][5] [12]),
        .I1(\slvo[6][hconfig][5] [12]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][5] [12]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][5] [12]),
        .O(\syncrregs.r[hrdatas][12]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][12]_i_27 
       (.I0(\slvo[3][hconfig][6] [12]),
        .I1(\slvo[2][hconfig][6] [12]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][6] [12]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][6] [12]),
        .O(\syncrregs.r[hrdatas][12]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][12]_i_28 
       (.I0(\slvo[7][hconfig][6] [12]),
        .I1(\slvo[6][hconfig][6] [12]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][6] [12]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][6] [12]),
        .O(\syncrregs.r[hrdatas][12]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][12]_i_29 
       (.I0(\slvo[3][hconfig][7] [12]),
        .I1(\slvo[2][hconfig][7] [12]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][7] [12]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][7] [12]),
        .O(\syncrregs.r[hrdatas][12]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \syncrregs.r[hrdatas][12]_i_3 
       (.I0(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I1(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I2(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I3(sel0[3]),
        .I4(sel0[5]),
        .I5(sel0[4]),
        .O(\syncrregs.r[hrdatas][12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][12]_i_30 
       (.I0(\slvo[7][hconfig][7] [12]),
        .I1(\slvo[6][hconfig][7] [12]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][7] [12]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][7] [12]),
        .O(\syncrregs.r[hrdatas][12]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][12]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][12]_i_7_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][12]_i_8_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I3(\syncrregs.r_reg[hrdatas][12]_i_9_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][2] ),
        .I5(\syncrregs.r_reg[hrdatas][12]_i_10_n_0 ),
        .O(\syncrregs.r[hrdatas][12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][13]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][13]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][13]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][13]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][13]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][13]_i_14 
       (.I0(\slvo[3][hconfig][6] [13]),
        .I1(\slvo[2][hconfig][6] [13]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][6] [13]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][6] [13]),
        .O(\syncrregs.r[hrdatas][13]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][13]_i_15 
       (.I0(\slvo[7][hconfig][6] [13]),
        .I1(\slvo[6][hconfig][6] [13]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][6] [13]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][6] [13]),
        .O(\syncrregs.r[hrdatas][13]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][13]_i_16 
       (.I0(\slvo[3][hconfig][7] [13]),
        .I1(\slvo[2][hconfig][7] [13]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][7] [13]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][7] [13]),
        .O(\syncrregs.r[hrdatas][13]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][13]_i_17 
       (.I0(\slvo[7][hconfig][7] [13]),
        .I1(\slvo[6][hconfig][7] [13]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][7] [13]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][7] [13]),
        .O(\syncrregs.r[hrdatas][13]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][13]_i_18 
       (.I0(\slvo[3][hconfig][4] [13]),
        .I1(\slvo[2][hconfig][4] [13]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][4] [13]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][4] [13]),
        .O(\syncrregs.r[hrdatas][13]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][13]_i_19 
       (.I0(\slvo[7][hconfig][4] [13]),
        .I1(\slvo[6][hconfig][4] [13]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][4] [13]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][4] [13]),
        .O(\syncrregs.r[hrdatas][13]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][13]_i_20 
       (.I0(\slvo[3][hconfig][5] [13]),
        .I1(\slvo[2][hconfig][5] [13]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][5] [13]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][5] [13]),
        .O(\syncrregs.r[hrdatas][13]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][13]_i_21 
       (.I0(\slvo[7][hconfig][5] [13]),
        .I1(\slvo[6][hconfig][5] [13]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][5] [13]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][5] [13]),
        .O(\syncrregs.r[hrdatas][13]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][13]_i_22 
       (.I0(\slvo[3][hconfig][2] [13]),
        .I1(\slvo[2][hconfig][2] [13]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][2] [13]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][2] [13]),
        .O(\syncrregs.r[hrdatas][13]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][13]_i_23 
       (.I0(\slvo[7][hconfig][2] [13]),
        .I1(\slvo[6][hconfig][2] [13]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][2] [13]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][2] [13]),
        .O(\syncrregs.r[hrdatas][13]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][13]_i_24 
       (.I0(\slvo[3][hconfig][3] [13]),
        .I1(\slvo[2][hconfig][3] [13]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][3] [13]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][3] [13]),
        .O(\syncrregs.r[hrdatas][13]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][13]_i_25 
       (.I0(\slvo[7][hconfig][3] [13]),
        .I1(\slvo[6][hconfig][3] [13]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][3] [13]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][3] [13]),
        .O(\syncrregs.r[hrdatas][13]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][13]_i_26 
       (.I0(\slvo[3][hconfig][0] [13]),
        .I1(\slvo[2][hconfig][0] [13]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][0] [13]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][0] [13]),
        .O(\syncrregs.r[hrdatas][13]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][13]_i_27 
       (.I0(\slvo[7][hconfig][0] [13]),
        .I1(\slvo[6][hconfig][0] [13]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][0] [13]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][0] [13]),
        .O(\syncrregs.r[hrdatas][13]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][13]_i_28 
       (.I0(\slvo[3][hconfig][1] [13]),
        .I1(\slvo[2][hconfig][1] [13]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][1] [13]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][1] [13]),
        .O(\syncrregs.r[hrdatas][13]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][13]_i_29 
       (.I0(\slvo[7][hconfig][1] [13]),
        .I1(\slvo[6][hconfig][1] [13]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][1] [13]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][1] [13]),
        .O(\syncrregs.r[hrdatas][13]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][14]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][14]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][14]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][14]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][14]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][14]_i_14 
       (.I0(\slvo[3][hconfig][6] [14]),
        .I1(\slvo[2][hconfig][6] [14]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][6] [14]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][6] [14]),
        .O(\syncrregs.r[hrdatas][14]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][14]_i_15 
       (.I0(\slvo[7][hconfig][6] [14]),
        .I1(\slvo[6][hconfig][6] [14]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][6] [14]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][6] [14]),
        .O(\syncrregs.r[hrdatas][14]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][14]_i_16 
       (.I0(\slvo[3][hconfig][7] [14]),
        .I1(\slvo[2][hconfig][7] [14]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][7] [14]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][7] [14]),
        .O(\syncrregs.r[hrdatas][14]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][14]_i_17 
       (.I0(\slvo[7][hconfig][7] [14]),
        .I1(\slvo[6][hconfig][7] [14]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][7] [14]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][7] [14]),
        .O(\syncrregs.r[hrdatas][14]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][14]_i_18 
       (.I0(\slvo[3][hconfig][4] [14]),
        .I1(\slvo[2][hconfig][4] [14]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][4] [14]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][4] [14]),
        .O(\syncrregs.r[hrdatas][14]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][14]_i_19 
       (.I0(\slvo[7][hconfig][4] [14]),
        .I1(\slvo[6][hconfig][4] [14]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][4] [14]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][4] [14]),
        .O(\syncrregs.r[hrdatas][14]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][14]_i_20 
       (.I0(\slvo[3][hconfig][5] [14]),
        .I1(\slvo[2][hconfig][5] [14]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][5] [14]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][5] [14]),
        .O(\syncrregs.r[hrdatas][14]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][14]_i_21 
       (.I0(\slvo[7][hconfig][5] [14]),
        .I1(\slvo[6][hconfig][5] [14]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][5] [14]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][5] [14]),
        .O(\syncrregs.r[hrdatas][14]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][14]_i_22 
       (.I0(\slvo[3][hconfig][2] [14]),
        .I1(\slvo[2][hconfig][2] [14]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][2] [14]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][2] [14]),
        .O(\syncrregs.r[hrdatas][14]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][14]_i_23 
       (.I0(\slvo[7][hconfig][2] [14]),
        .I1(\slvo[6][hconfig][2] [14]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][2] [14]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][2] [14]),
        .O(\syncrregs.r[hrdatas][14]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][14]_i_24 
       (.I0(\slvo[3][hconfig][3] [14]),
        .I1(\slvo[2][hconfig][3] [14]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][3] [14]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][3] [14]),
        .O(\syncrregs.r[hrdatas][14]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][14]_i_25 
       (.I0(\slvo[7][hconfig][3] [14]),
        .I1(\slvo[6][hconfig][3] [14]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][3] [14]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][3] [14]),
        .O(\syncrregs.r[hrdatas][14]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][14]_i_26 
       (.I0(\slvo[3][hconfig][0] [14]),
        .I1(\slvo[2][hconfig][0] [14]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][0] [14]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][0] [14]),
        .O(\syncrregs.r[hrdatas][14]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][14]_i_27 
       (.I0(\slvo[7][hconfig][0] [14]),
        .I1(\slvo[6][hconfig][0] [14]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][0] [14]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][0] [14]),
        .O(\syncrregs.r[hrdatas][14]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][14]_i_28 
       (.I0(\slvo[3][hconfig][1] [14]),
        .I1(\slvo[2][hconfig][1] [14]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][1] [14]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][1] [14]),
        .O(\syncrregs.r[hrdatas][14]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][14]_i_29 
       (.I0(\slvo[7][hconfig][1] [14]),
        .I1(\slvo[6][hconfig][1] [14]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][1] [14]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][1] [14]),
        .O(\syncrregs.r[hrdatas][14]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][15]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][15]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][15]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][15]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][15]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][15]_i_14 
       (.I0(\slvo[3][hconfig][6] [15]),
        .I1(\slvo[2][hconfig][6] [15]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][6] [15]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][6] [15]),
        .O(\syncrregs.r[hrdatas][15]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][15]_i_15 
       (.I0(\slvo[7][hconfig][6] [15]),
        .I1(\slvo[6][hconfig][6] [15]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][6] [15]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][6] [15]),
        .O(\syncrregs.r[hrdatas][15]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][15]_i_16 
       (.I0(\slvo[3][hconfig][7] [15]),
        .I1(\slvo[2][hconfig][7] [15]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][7] [15]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][7] [15]),
        .O(\syncrregs.r[hrdatas][15]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][15]_i_17 
       (.I0(\slvo[7][hconfig][7] [15]),
        .I1(\slvo[6][hconfig][7] [15]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][7] [15]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][7] [15]),
        .O(\syncrregs.r[hrdatas][15]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][15]_i_18 
       (.I0(\slvo[3][hconfig][4] [15]),
        .I1(\slvo[2][hconfig][4] [15]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][4] [15]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][4] [15]),
        .O(\syncrregs.r[hrdatas][15]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][15]_i_19 
       (.I0(\slvo[7][hconfig][4] [15]),
        .I1(\slvo[6][hconfig][4] [15]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][4] [15]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][4] [15]),
        .O(\syncrregs.r[hrdatas][15]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][15]_i_20 
       (.I0(\slvo[3][hconfig][5] [15]),
        .I1(\slvo[2][hconfig][5] [15]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][5] [15]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][5] [15]),
        .O(\syncrregs.r[hrdatas][15]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][15]_i_21 
       (.I0(\slvo[7][hconfig][5] [15]),
        .I1(\slvo[6][hconfig][5] [15]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][5] [15]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][5] [15]),
        .O(\syncrregs.r[hrdatas][15]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][15]_i_22 
       (.I0(\slvo[3][hconfig][2] [15]),
        .I1(\slvo[2][hconfig][2] [15]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][2] [15]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][2] [15]),
        .O(\syncrregs.r[hrdatas][15]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][15]_i_23 
       (.I0(\slvo[7][hconfig][2] [15]),
        .I1(\slvo[6][hconfig][2] [15]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][2] [15]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][2] [15]),
        .O(\syncrregs.r[hrdatas][15]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][15]_i_24 
       (.I0(\slvo[3][hconfig][3] [15]),
        .I1(\slvo[2][hconfig][3] [15]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][3] [15]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][3] [15]),
        .O(\syncrregs.r[hrdatas][15]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][15]_i_25 
       (.I0(\slvo[7][hconfig][3] [15]),
        .I1(\slvo[6][hconfig][3] [15]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][3] [15]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][3] [15]),
        .O(\syncrregs.r[hrdatas][15]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][15]_i_26 
       (.I0(\slvo[3][hconfig][0] [15]),
        .I1(\slvo[2][hconfig][0] [15]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][0] [15]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][0] [15]),
        .O(\syncrregs.r[hrdatas][15]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][15]_i_27 
       (.I0(\slvo[7][hconfig][0] [15]),
        .I1(\slvo[6][hconfig][0] [15]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][0] [15]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][0] [15]),
        .O(\syncrregs.r[hrdatas][15]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][15]_i_28 
       (.I0(\slvo[3][hconfig][1] [15]),
        .I1(\slvo[2][hconfig][1] [15]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][1] [15]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][1] [15]),
        .O(\syncrregs.r[hrdatas][15]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][15]_i_29 
       (.I0(\slvo[7][hconfig][1] [15]),
        .I1(\slvo[6][hconfig][1] [15]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][1] [15]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][1] [15]),
        .O(\syncrregs.r[hrdatas][15]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][16]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][16]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][16]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][16]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][16]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][16]_i_14 
       (.I0(\slvo[3][hconfig][6] [16]),
        .I1(\slvo[2][hconfig][6] [16]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][6] [16]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][6] [16]),
        .O(\syncrregs.r[hrdatas][16]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][16]_i_15 
       (.I0(\slvo[7][hconfig][6] [16]),
        .I1(\slvo[6][hconfig][6] [16]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][6] [16]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][6] [16]),
        .O(\syncrregs.r[hrdatas][16]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][16]_i_16 
       (.I0(\slvo[3][hconfig][7] [16]),
        .I1(\slvo[2][hconfig][7] [16]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][7] [16]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][7] [16]),
        .O(\syncrregs.r[hrdatas][16]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][16]_i_17 
       (.I0(\slvo[7][hconfig][7] [16]),
        .I1(\slvo[6][hconfig][7] [16]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][7] [16]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][7] [16]),
        .O(\syncrregs.r[hrdatas][16]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][16]_i_18 
       (.I0(\slvo[3][hconfig][4] [16]),
        .I1(\slvo[2][hconfig][4] [16]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][4] [16]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][4] [16]),
        .O(\syncrregs.r[hrdatas][16]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][16]_i_19 
       (.I0(\slvo[7][hconfig][4] [16]),
        .I1(\slvo[6][hconfig][4] [16]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][4] [16]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][4] [16]),
        .O(\syncrregs.r[hrdatas][16]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][16]_i_20 
       (.I0(\slvo[3][hconfig][5] [16]),
        .I1(\slvo[2][hconfig][5] [16]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][5] [16]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][5] [16]),
        .O(\syncrregs.r[hrdatas][16]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][16]_i_21 
       (.I0(\slvo[7][hconfig][5] [16]),
        .I1(\slvo[6][hconfig][5] [16]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][5] [16]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][5] [16]),
        .O(\syncrregs.r[hrdatas][16]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][16]_i_22 
       (.I0(\slvo[3][hconfig][2] [16]),
        .I1(\slvo[2][hconfig][2] [16]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][2] [16]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][2] [16]),
        .O(\syncrregs.r[hrdatas][16]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][16]_i_23 
       (.I0(\slvo[7][hconfig][2] [16]),
        .I1(\slvo[6][hconfig][2] [16]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][2] [16]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][2] [16]),
        .O(\syncrregs.r[hrdatas][16]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][16]_i_24 
       (.I0(\slvo[3][hconfig][3] [16]),
        .I1(\slvo[2][hconfig][3] [16]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][3] [16]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][3] [16]),
        .O(\syncrregs.r[hrdatas][16]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][16]_i_25 
       (.I0(\slvo[7][hconfig][3] [16]),
        .I1(\slvo[6][hconfig][3] [16]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][3] [16]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][3] [16]),
        .O(\syncrregs.r[hrdatas][16]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][16]_i_26 
       (.I0(\slvo[3][hconfig][0] [16]),
        .I1(\slvo[2][hconfig][0] [16]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][0] [16]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][0] [16]),
        .O(\syncrregs.r[hrdatas][16]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][16]_i_27 
       (.I0(\slvo[7][hconfig][0] [16]),
        .I1(\slvo[6][hconfig][0] [16]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][0] [16]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][0] [16]),
        .O(\syncrregs.r[hrdatas][16]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][16]_i_28 
       (.I0(\slvo[3][hconfig][1] [16]),
        .I1(\slvo[2][hconfig][1] [16]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][1] [16]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][1] [16]),
        .O(\syncrregs.r[hrdatas][16]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][16]_i_29 
       (.I0(\slvo[7][hconfig][1] [16]),
        .I1(\slvo[6][hconfig][1] [16]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][1] [16]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][1] [16]),
        .O(\syncrregs.r[hrdatas][16]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][17]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][17]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][17]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][17]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][17]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][17]_i_14 
       (.I0(\slvo[3][hconfig][6] [17]),
        .I1(\slvo[2][hconfig][6] [17]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][6] [17]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][6] [17]),
        .O(\syncrregs.r[hrdatas][17]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][17]_i_15 
       (.I0(\slvo[7][hconfig][6] [17]),
        .I1(\slvo[6][hconfig][6] [17]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][6] [17]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][6] [17]),
        .O(\syncrregs.r[hrdatas][17]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][17]_i_16 
       (.I0(\slvo[3][hconfig][7] [17]),
        .I1(\slvo[2][hconfig][7] [17]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][7] [17]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][7] [17]),
        .O(\syncrregs.r[hrdatas][17]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][17]_i_17 
       (.I0(\slvo[7][hconfig][7] [17]),
        .I1(\slvo[6][hconfig][7] [17]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][7] [17]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][7] [17]),
        .O(\syncrregs.r[hrdatas][17]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][17]_i_18 
       (.I0(\slvo[3][hconfig][4] [17]),
        .I1(\slvo[2][hconfig][4] [17]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][4] [17]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][4] [17]),
        .O(\syncrregs.r[hrdatas][17]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][17]_i_19 
       (.I0(\slvo[7][hconfig][4] [17]),
        .I1(\slvo[6][hconfig][4] [17]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][4] [17]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][4] [17]),
        .O(\syncrregs.r[hrdatas][17]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][17]_i_20 
       (.I0(\slvo[3][hconfig][5] [17]),
        .I1(\slvo[2][hconfig][5] [17]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][5] [17]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][5] [17]),
        .O(\syncrregs.r[hrdatas][17]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][17]_i_21 
       (.I0(\slvo[7][hconfig][5] [17]),
        .I1(\slvo[6][hconfig][5] [17]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][5] [17]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][5] [17]),
        .O(\syncrregs.r[hrdatas][17]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][17]_i_22 
       (.I0(\slvo[3][hconfig][2] [17]),
        .I1(\slvo[2][hconfig][2] [17]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][2] [17]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][2] [17]),
        .O(\syncrregs.r[hrdatas][17]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][17]_i_23 
       (.I0(\slvo[7][hconfig][2] [17]),
        .I1(\slvo[6][hconfig][2] [17]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][2] [17]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][2] [17]),
        .O(\syncrregs.r[hrdatas][17]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][17]_i_24 
       (.I0(\slvo[3][hconfig][3] [17]),
        .I1(\slvo[2][hconfig][3] [17]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][3] [17]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][3] [17]),
        .O(\syncrregs.r[hrdatas][17]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][17]_i_25 
       (.I0(\slvo[7][hconfig][3] [17]),
        .I1(\slvo[6][hconfig][3] [17]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][3] [17]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][3] [17]),
        .O(\syncrregs.r[hrdatas][17]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][17]_i_26 
       (.I0(\slvo[3][hconfig][0] [17]),
        .I1(\slvo[2][hconfig][0] [17]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][0] [17]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][0] [17]),
        .O(\syncrregs.r[hrdatas][17]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][17]_i_27 
       (.I0(\slvo[7][hconfig][0] [17]),
        .I1(\slvo[6][hconfig][0] [17]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][0] [17]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][0] [17]),
        .O(\syncrregs.r[hrdatas][17]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][17]_i_28 
       (.I0(\slvo[3][hconfig][1] [17]),
        .I1(\slvo[2][hconfig][1] [17]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[1][hconfig][1] [17]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[0][hconfig][1] [17]),
        .O(\syncrregs.r[hrdatas][17]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][17]_i_29 
       (.I0(\slvo[7][hconfig][1] [17]),
        .I1(\slvo[6][hconfig][1] [17]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .I3(\slvo[5][hconfig][1] [17]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .I5(\slvo[4][hconfig][1] [17]),
        .O(\syncrregs.r[hrdatas][17]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][18]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][18]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][18]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][18]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][18]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][18]_i_14 
       (.I0(\slvo[3][hconfig][6] [18]),
        .I1(\slvo[2][hconfig][6] [18]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][6] [18]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][6] [18]),
        .O(\syncrregs.r[hrdatas][18]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][18]_i_15 
       (.I0(\slvo[7][hconfig][6] [18]),
        .I1(\slvo[6][hconfig][6] [18]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][6] [18]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][6] [18]),
        .O(\syncrregs.r[hrdatas][18]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][18]_i_16 
       (.I0(\slvo[3][hconfig][7] [18]),
        .I1(\slvo[2][hconfig][7] [18]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][7] [18]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][7] [18]),
        .O(\syncrregs.r[hrdatas][18]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][18]_i_17 
       (.I0(\slvo[7][hconfig][7] [18]),
        .I1(\slvo[6][hconfig][7] [18]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][7] [18]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][7] [18]),
        .O(\syncrregs.r[hrdatas][18]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][18]_i_18 
       (.I0(\slvo[3][hconfig][4] [18]),
        .I1(\slvo[2][hconfig][4] [18]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][4] [18]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][4] [18]),
        .O(\syncrregs.r[hrdatas][18]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][18]_i_19 
       (.I0(\slvo[7][hconfig][4] [18]),
        .I1(\slvo[6][hconfig][4] [18]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][4] [18]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][4] [18]),
        .O(\syncrregs.r[hrdatas][18]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][18]_i_20 
       (.I0(\slvo[3][hconfig][5] [18]),
        .I1(\slvo[2][hconfig][5] [18]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][5] [18]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][5] [18]),
        .O(\syncrregs.r[hrdatas][18]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][18]_i_21 
       (.I0(\slvo[7][hconfig][5] [18]),
        .I1(\slvo[6][hconfig][5] [18]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][5] [18]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][5] [18]),
        .O(\syncrregs.r[hrdatas][18]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][18]_i_22 
       (.I0(\slvo[3][hconfig][2] [18]),
        .I1(\slvo[2][hconfig][2] [18]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][2] [18]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][2] [18]),
        .O(\syncrregs.r[hrdatas][18]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][18]_i_23 
       (.I0(\slvo[7][hconfig][2] [18]),
        .I1(\slvo[6][hconfig][2] [18]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][2] [18]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][2] [18]),
        .O(\syncrregs.r[hrdatas][18]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][18]_i_24 
       (.I0(\slvo[3][hconfig][3] [18]),
        .I1(\slvo[2][hconfig][3] [18]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][3] [18]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][3] [18]),
        .O(\syncrregs.r[hrdatas][18]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][18]_i_25 
       (.I0(\slvo[7][hconfig][3] [18]),
        .I1(\slvo[6][hconfig][3] [18]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][3] [18]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][3] [18]),
        .O(\syncrregs.r[hrdatas][18]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][18]_i_26 
       (.I0(\slvo[3][hconfig][0] [18]),
        .I1(\slvo[2][hconfig][0] [18]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][0] [18]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][0] [18]),
        .O(\syncrregs.r[hrdatas][18]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][18]_i_27 
       (.I0(\slvo[7][hconfig][0] [18]),
        .I1(\slvo[6][hconfig][0] [18]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][0] [18]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][0] [18]),
        .O(\syncrregs.r[hrdatas][18]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][18]_i_28 
       (.I0(\slvo[3][hconfig][1] [18]),
        .I1(\slvo[2][hconfig][1] [18]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][1] [18]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][1] [18]),
        .O(\syncrregs.r[hrdatas][18]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][18]_i_29 
       (.I0(\slvo[7][hconfig][1] [18]),
        .I1(\slvo[6][hconfig][1] [18]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][1] [18]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][1] [18]),
        .O(\syncrregs.r[hrdatas][18]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][19]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][19]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][19]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][19]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][19]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][19]_i_14 
       (.I0(\slvo[3][hconfig][6] [19]),
        .I1(\slvo[2][hconfig][6] [19]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][6] [19]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][6] [19]),
        .O(\syncrregs.r[hrdatas][19]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][19]_i_15 
       (.I0(\slvo[7][hconfig][6] [19]),
        .I1(\slvo[6][hconfig][6] [19]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][6] [19]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][6] [19]),
        .O(\syncrregs.r[hrdatas][19]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][19]_i_16 
       (.I0(\slvo[3][hconfig][7] [19]),
        .I1(\slvo[2][hconfig][7] [19]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][7] [19]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][7] [19]),
        .O(\syncrregs.r[hrdatas][19]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][19]_i_17 
       (.I0(\slvo[7][hconfig][7] [19]),
        .I1(\slvo[6][hconfig][7] [19]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][7] [19]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][7] [19]),
        .O(\syncrregs.r[hrdatas][19]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][19]_i_18 
       (.I0(\slvo[3][hconfig][4] [19]),
        .I1(\slvo[2][hconfig][4] [19]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][4] [19]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][4] [19]),
        .O(\syncrregs.r[hrdatas][19]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][19]_i_19 
       (.I0(\slvo[7][hconfig][4] [19]),
        .I1(\slvo[6][hconfig][4] [19]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][4] [19]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][4] [19]),
        .O(\syncrregs.r[hrdatas][19]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][19]_i_20 
       (.I0(\slvo[3][hconfig][5] [19]),
        .I1(\slvo[2][hconfig][5] [19]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][5] [19]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][5] [19]),
        .O(\syncrregs.r[hrdatas][19]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][19]_i_21 
       (.I0(\slvo[7][hconfig][5] [19]),
        .I1(\slvo[6][hconfig][5] [19]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][5] [19]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][5] [19]),
        .O(\syncrregs.r[hrdatas][19]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][19]_i_22 
       (.I0(\slvo[3][hconfig][2] [19]),
        .I1(\slvo[2][hconfig][2] [19]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][2] [19]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][2] [19]),
        .O(\syncrregs.r[hrdatas][19]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][19]_i_23 
       (.I0(\slvo[7][hconfig][2] [19]),
        .I1(\slvo[6][hconfig][2] [19]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][2] [19]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][2] [19]),
        .O(\syncrregs.r[hrdatas][19]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][19]_i_24 
       (.I0(\slvo[3][hconfig][3] [19]),
        .I1(\slvo[2][hconfig][3] [19]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][3] [19]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][3] [19]),
        .O(\syncrregs.r[hrdatas][19]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][19]_i_25 
       (.I0(\slvo[7][hconfig][3] [19]),
        .I1(\slvo[6][hconfig][3] [19]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][3] [19]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][3] [19]),
        .O(\syncrregs.r[hrdatas][19]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][19]_i_26 
       (.I0(\slvo[3][hconfig][0] [19]),
        .I1(\slvo[2][hconfig][0] [19]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][0] [19]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][0] [19]),
        .O(\syncrregs.r[hrdatas][19]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][19]_i_27 
       (.I0(\slvo[7][hconfig][0] [19]),
        .I1(\slvo[6][hconfig][0] [19]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][0] [19]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][0] [19]),
        .O(\syncrregs.r[hrdatas][19]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][19]_i_28 
       (.I0(\slvo[3][hconfig][1] [19]),
        .I1(\slvo[2][hconfig][1] [19]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][1] [19]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][1] [19]),
        .O(\syncrregs.r[hrdatas][19]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][19]_i_29 
       (.I0(\slvo[7][hconfig][1] [19]),
        .I1(\slvo[6][hconfig][1] [19]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][1] [19]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][1] [19]),
        .O(\syncrregs.r[hrdatas][19]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEE222E200000000)) 
    \syncrregs.r[hrdatas][1]_i_1 
       (.I0(\syncrregs.r[hrdatas][1]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I2(\syncrregs.r_reg[hrdatas][1]_i_3_n_0 ),
        .I3(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I4(\syncrregs.r_reg[hrdatas][1]_i_4_n_0 ),
        .I5(p_179_out),
        .O(\syncrregs.r[hrdatas][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][1]_i_13 
       (.I0(\slvo[3][hconfig][3] [1]),
        .I1(\slvo[2][hconfig][3] [1]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][3] [1]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][3] [1]),
        .O(\syncrregs.r[hrdatas][1]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][1]_i_14 
       (.I0(\slvo[7][hconfig][3] [1]),
        .I1(\slvo[6][hconfig][3] [1]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][3] [1]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][3] [1]),
        .O(\syncrregs.r[hrdatas][1]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][1]_i_15 
       (.I0(\slvo[3][hconfig][2] [1]),
        .I1(\slvo[2][hconfig][2] [1]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][2] [1]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][2] [1]),
        .O(\syncrregs.r[hrdatas][1]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][1]_i_16 
       (.I0(\slvo[7][hconfig][2] [1]),
        .I1(\slvo[6][hconfig][2] [1]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][2] [1]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][2] [1]),
        .O(\syncrregs.r[hrdatas][1]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][1]_i_17 
       (.I0(\slvo[3][hconfig][1] [1]),
        .I1(\slvo[2][hconfig][1] [1]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][1] [1]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][1] [1]),
        .O(\syncrregs.r[hrdatas][1]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][1]_i_18 
       (.I0(\slvo[7][hconfig][1] [1]),
        .I1(\slvo[6][hconfig][1] [1]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][1] [1]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][1] [1]),
        .O(\syncrregs.r[hrdatas][1]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][1]_i_19 
       (.I0(\slvo[3][hconfig][0] [1]),
        .I1(\slvo[2][hconfig][0] [1]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][0] [1]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][0] [1]),
        .O(\syncrregs.r[hrdatas][1]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][1]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][1]_i_5_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][1]_i_6_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I3(\syncrregs.r_reg[hrdatas][1]_i_7_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][2] ),
        .I5(\syncrregs.r_reg[hrdatas][1]_i_8_n_0 ),
        .O(\syncrregs.r[hrdatas][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][1]_i_20 
       (.I0(\slvo[7][hconfig][0] [1]),
        .I1(\slvo[6][hconfig][0] [1]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][0] [1]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][0] [1]),
        .O(\syncrregs.r[hrdatas][1]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][1]_i_21 
       (.I0(\slvo[3][hconfig][4] [1]),
        .I1(\slvo[2][hconfig][4] [1]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][4] [1]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][4] [1]),
        .O(\syncrregs.r[hrdatas][1]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][1]_i_22 
       (.I0(\slvo[7][hconfig][4] [1]),
        .I1(\slvo[6][hconfig][4] [1]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][4] [1]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][4] [1]),
        .O(\syncrregs.r[hrdatas][1]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][1]_i_23 
       (.I0(\slvo[3][hconfig][5] [1]),
        .I1(\slvo[2][hconfig][5] [1]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][5] [1]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][5] [1]),
        .O(\syncrregs.r[hrdatas][1]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][1]_i_24 
       (.I0(\slvo[7][hconfig][5] [1]),
        .I1(\slvo[6][hconfig][5] [1]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][5] [1]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][5] [1]),
        .O(\syncrregs.r[hrdatas][1]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][1]_i_25 
       (.I0(\slvo[3][hconfig][6] [1]),
        .I1(\slvo[2][hconfig][6] [1]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][6] [1]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][6] [1]),
        .O(\syncrregs.r[hrdatas][1]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][1]_i_26 
       (.I0(\slvo[7][hconfig][6] [1]),
        .I1(\slvo[6][hconfig][6] [1]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][6] [1]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][6] [1]),
        .O(\syncrregs.r[hrdatas][1]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][1]_i_27 
       (.I0(\slvo[3][hconfig][7] [1]),
        .I1(\slvo[2][hconfig][7] [1]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][7] [1]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][7] [1]),
        .O(\syncrregs.r[hrdatas][1]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][1]_i_28 
       (.I0(\slvo[7][hconfig][7] [1]),
        .I1(\slvo[6][hconfig][7] [1]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][7] [1]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][7] [1]),
        .O(\syncrregs.r[hrdatas][1]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][20]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][20]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][20]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][20]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][20]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][20]_i_14 
       (.I0(\slvo[3][hconfig][6] [20]),
        .I1(\slvo[2][hconfig][6] [20]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][6] [20]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][6] [20]),
        .O(\syncrregs.r[hrdatas][20]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][20]_i_15 
       (.I0(\slvo[7][hconfig][6] [20]),
        .I1(\slvo[6][hconfig][6] [20]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][6] [20]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][6] [20]),
        .O(\syncrregs.r[hrdatas][20]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][20]_i_16 
       (.I0(\slvo[3][hconfig][7] [20]),
        .I1(\slvo[2][hconfig][7] [20]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][7] [20]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][7] [20]),
        .O(\syncrregs.r[hrdatas][20]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][20]_i_17 
       (.I0(\slvo[7][hconfig][7] [20]),
        .I1(\slvo[6][hconfig][7] [20]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][7] [20]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][7] [20]),
        .O(\syncrregs.r[hrdatas][20]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][20]_i_18 
       (.I0(\slvo[3][hconfig][4] [20]),
        .I1(\slvo[2][hconfig][4] [20]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][4] [20]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][4] [20]),
        .O(\syncrregs.r[hrdatas][20]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][20]_i_19 
       (.I0(\slvo[7][hconfig][4] [20]),
        .I1(\slvo[6][hconfig][4] [20]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][4] [20]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][4] [20]),
        .O(\syncrregs.r[hrdatas][20]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][20]_i_20 
       (.I0(\slvo[3][hconfig][5] [20]),
        .I1(\slvo[2][hconfig][5] [20]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][5] [20]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][5] [20]),
        .O(\syncrregs.r[hrdatas][20]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][20]_i_21 
       (.I0(\slvo[7][hconfig][5] [20]),
        .I1(\slvo[6][hconfig][5] [20]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][5] [20]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][5] [20]),
        .O(\syncrregs.r[hrdatas][20]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][20]_i_22 
       (.I0(\slvo[3][hconfig][2] [20]),
        .I1(\slvo[2][hconfig][2] [20]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][2] [20]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][2] [20]),
        .O(\syncrregs.r[hrdatas][20]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][20]_i_23 
       (.I0(\slvo[7][hconfig][2] [20]),
        .I1(\slvo[6][hconfig][2] [20]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][2] [20]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][2] [20]),
        .O(\syncrregs.r[hrdatas][20]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][20]_i_24 
       (.I0(\slvo[3][hconfig][3] [20]),
        .I1(\slvo[2][hconfig][3] [20]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][3] [20]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][3] [20]),
        .O(\syncrregs.r[hrdatas][20]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][20]_i_25 
       (.I0(\slvo[7][hconfig][3] [20]),
        .I1(\slvo[6][hconfig][3] [20]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][3] [20]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][3] [20]),
        .O(\syncrregs.r[hrdatas][20]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][20]_i_26 
       (.I0(\slvo[3][hconfig][0] [20]),
        .I1(\slvo[2][hconfig][0] [20]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][0] [20]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][0] [20]),
        .O(\syncrregs.r[hrdatas][20]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][20]_i_27 
       (.I0(\slvo[7][hconfig][0] [20]),
        .I1(\slvo[6][hconfig][0] [20]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][0] [20]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][0] [20]),
        .O(\syncrregs.r[hrdatas][20]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][20]_i_28 
       (.I0(\slvo[3][hconfig][1] [20]),
        .I1(\slvo[2][hconfig][1] [20]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][1] [20]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][1] [20]),
        .O(\syncrregs.r[hrdatas][20]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][20]_i_29 
       (.I0(\slvo[7][hconfig][1] [20]),
        .I1(\slvo[6][hconfig][1] [20]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][1] [20]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][1] [20]),
        .O(\syncrregs.r[hrdatas][20]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][21]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][21]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][21]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][21]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][21]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][21]_i_14 
       (.I0(\slvo[3][hconfig][6] [21]),
        .I1(\slvo[2][hconfig][6] [21]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][6] [21]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][6] [21]),
        .O(\syncrregs.r[hrdatas][21]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][21]_i_15 
       (.I0(\slvo[7][hconfig][6] [21]),
        .I1(\slvo[6][hconfig][6] [21]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][6] [21]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][6] [21]),
        .O(\syncrregs.r[hrdatas][21]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][21]_i_16 
       (.I0(\slvo[3][hconfig][7] [21]),
        .I1(\slvo[2][hconfig][7] [21]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][7] [21]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][7] [21]),
        .O(\syncrregs.r[hrdatas][21]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][21]_i_17 
       (.I0(\slvo[7][hconfig][7] [21]),
        .I1(\slvo[6][hconfig][7] [21]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][7] [21]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][7] [21]),
        .O(\syncrregs.r[hrdatas][21]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][21]_i_18 
       (.I0(\slvo[3][hconfig][4] [21]),
        .I1(\slvo[2][hconfig][4] [21]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][4] [21]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][4] [21]),
        .O(\syncrregs.r[hrdatas][21]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][21]_i_19 
       (.I0(\slvo[7][hconfig][4] [21]),
        .I1(\slvo[6][hconfig][4] [21]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][4] [21]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][4] [21]),
        .O(\syncrregs.r[hrdatas][21]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][21]_i_20 
       (.I0(\slvo[3][hconfig][5] [21]),
        .I1(\slvo[2][hconfig][5] [21]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][5] [21]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][5] [21]),
        .O(\syncrregs.r[hrdatas][21]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][21]_i_21 
       (.I0(\slvo[7][hconfig][5] [21]),
        .I1(\slvo[6][hconfig][5] [21]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][5] [21]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][5] [21]),
        .O(\syncrregs.r[hrdatas][21]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][21]_i_22 
       (.I0(\slvo[3][hconfig][2] [21]),
        .I1(\slvo[2][hconfig][2] [21]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][2] [21]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][2] [21]),
        .O(\syncrregs.r[hrdatas][21]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][21]_i_23 
       (.I0(\slvo[7][hconfig][2] [21]),
        .I1(\slvo[6][hconfig][2] [21]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][2] [21]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][2] [21]),
        .O(\syncrregs.r[hrdatas][21]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][21]_i_24 
       (.I0(\slvo[3][hconfig][3] [21]),
        .I1(\slvo[2][hconfig][3] [21]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][3] [21]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][3] [21]),
        .O(\syncrregs.r[hrdatas][21]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][21]_i_25 
       (.I0(\slvo[7][hconfig][3] [21]),
        .I1(\slvo[6][hconfig][3] [21]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][3] [21]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][3] [21]),
        .O(\syncrregs.r[hrdatas][21]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][21]_i_26 
       (.I0(\slvo[3][hconfig][0] [21]),
        .I1(\slvo[2][hconfig][0] [21]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][0] [21]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][0] [21]),
        .O(\syncrregs.r[hrdatas][21]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][21]_i_27 
       (.I0(\slvo[7][hconfig][0] [21]),
        .I1(\slvo[6][hconfig][0] [21]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][0] [21]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][0] [21]),
        .O(\syncrregs.r[hrdatas][21]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][21]_i_28 
       (.I0(\slvo[3][hconfig][1] [21]),
        .I1(\slvo[2][hconfig][1] [21]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][1] [21]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][1] [21]),
        .O(\syncrregs.r[hrdatas][21]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][21]_i_29 
       (.I0(\slvo[7][hconfig][1] [21]),
        .I1(\slvo[6][hconfig][1] [21]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][1] [21]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][1] [21]),
        .O(\syncrregs.r[hrdatas][21]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][22]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][22]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][22]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][22]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][22]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][22]_i_14 
       (.I0(\slvo[3][hconfig][6] [22]),
        .I1(\slvo[2][hconfig][6] [22]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][6] [22]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][6] [22]),
        .O(\syncrregs.r[hrdatas][22]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][22]_i_15 
       (.I0(\slvo[7][hconfig][6] [22]),
        .I1(\slvo[6][hconfig][6] [22]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][6] [22]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][6] [22]),
        .O(\syncrregs.r[hrdatas][22]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][22]_i_16 
       (.I0(\slvo[3][hconfig][7] [22]),
        .I1(\slvo[2][hconfig][7] [22]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][7] [22]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][7] [22]),
        .O(\syncrregs.r[hrdatas][22]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][22]_i_17 
       (.I0(\slvo[7][hconfig][7] [22]),
        .I1(\slvo[6][hconfig][7] [22]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][7] [22]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][7] [22]),
        .O(\syncrregs.r[hrdatas][22]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][22]_i_18 
       (.I0(\slvo[3][hconfig][4] [22]),
        .I1(\slvo[2][hconfig][4] [22]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][4] [22]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][4] [22]),
        .O(\syncrregs.r[hrdatas][22]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][22]_i_19 
       (.I0(\slvo[7][hconfig][4] [22]),
        .I1(\slvo[6][hconfig][4] [22]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][4] [22]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][4] [22]),
        .O(\syncrregs.r[hrdatas][22]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][22]_i_20 
       (.I0(\slvo[3][hconfig][5] [22]),
        .I1(\slvo[2][hconfig][5] [22]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][5] [22]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][5] [22]),
        .O(\syncrregs.r[hrdatas][22]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][22]_i_21 
       (.I0(\slvo[7][hconfig][5] [22]),
        .I1(\slvo[6][hconfig][5] [22]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][5] [22]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][5] [22]),
        .O(\syncrregs.r[hrdatas][22]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][22]_i_22 
       (.I0(\slvo[3][hconfig][2] [22]),
        .I1(\slvo[2][hconfig][2] [22]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][2] [22]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][2] [22]),
        .O(\syncrregs.r[hrdatas][22]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][22]_i_23 
       (.I0(\slvo[7][hconfig][2] [22]),
        .I1(\slvo[6][hconfig][2] [22]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][2] [22]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][2] [22]),
        .O(\syncrregs.r[hrdatas][22]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][22]_i_24 
       (.I0(\slvo[3][hconfig][3] [22]),
        .I1(\slvo[2][hconfig][3] [22]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][3] [22]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][3] [22]),
        .O(\syncrregs.r[hrdatas][22]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][22]_i_25 
       (.I0(\slvo[7][hconfig][3] [22]),
        .I1(\slvo[6][hconfig][3] [22]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][3] [22]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][3] [22]),
        .O(\syncrregs.r[hrdatas][22]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][22]_i_26 
       (.I0(\slvo[3][hconfig][0] [22]),
        .I1(\slvo[2][hconfig][0] [22]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][0] [22]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][0] [22]),
        .O(\syncrregs.r[hrdatas][22]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][22]_i_27 
       (.I0(\slvo[7][hconfig][0] [22]),
        .I1(\slvo[6][hconfig][0] [22]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][0] [22]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][0] [22]),
        .O(\syncrregs.r[hrdatas][22]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][22]_i_28 
       (.I0(\slvo[3][hconfig][1] [22]),
        .I1(\slvo[2][hconfig][1] [22]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][1] [22]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][1] [22]),
        .O(\syncrregs.r[hrdatas][22]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][22]_i_29 
       (.I0(\slvo[7][hconfig][1] [22]),
        .I1(\slvo[6][hconfig][1] [22]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][1] [22]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][1] [22]),
        .O(\syncrregs.r[hrdatas][22]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][23]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][23]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][23]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][23]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][23]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][23]_i_14 
       (.I0(\slvo[3][hconfig][6] [23]),
        .I1(\slvo[2][hconfig][6] [23]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][6] [23]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][6] [23]),
        .O(\syncrregs.r[hrdatas][23]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][23]_i_15 
       (.I0(\slvo[7][hconfig][6] [23]),
        .I1(\slvo[6][hconfig][6] [23]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][6] [23]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][6] [23]),
        .O(\syncrregs.r[hrdatas][23]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][23]_i_16 
       (.I0(\slvo[3][hconfig][7] [23]),
        .I1(\slvo[2][hconfig][7] [23]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][7] [23]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][7] [23]),
        .O(\syncrregs.r[hrdatas][23]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][23]_i_17 
       (.I0(\slvo[7][hconfig][7] [23]),
        .I1(\slvo[6][hconfig][7] [23]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][7] [23]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][7] [23]),
        .O(\syncrregs.r[hrdatas][23]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][23]_i_18 
       (.I0(\slvo[3][hconfig][4] [23]),
        .I1(\slvo[2][hconfig][4] [23]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][4] [23]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][4] [23]),
        .O(\syncrregs.r[hrdatas][23]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][23]_i_19 
       (.I0(\slvo[7][hconfig][4] [23]),
        .I1(\slvo[6][hconfig][4] [23]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][4] [23]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][4] [23]),
        .O(\syncrregs.r[hrdatas][23]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][23]_i_20 
       (.I0(\slvo[3][hconfig][5] [23]),
        .I1(\slvo[2][hconfig][5] [23]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][5] [23]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][5] [23]),
        .O(\syncrregs.r[hrdatas][23]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][23]_i_21 
       (.I0(\slvo[7][hconfig][5] [23]),
        .I1(\slvo[6][hconfig][5] [23]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][5] [23]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][5] [23]),
        .O(\syncrregs.r[hrdatas][23]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][23]_i_22 
       (.I0(\slvo[3][hconfig][2] [23]),
        .I1(\slvo[2][hconfig][2] [23]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][2] [23]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][2] [23]),
        .O(\syncrregs.r[hrdatas][23]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][23]_i_23 
       (.I0(\slvo[7][hconfig][2] [23]),
        .I1(\slvo[6][hconfig][2] [23]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][2] [23]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][2] [23]),
        .O(\syncrregs.r[hrdatas][23]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][23]_i_24 
       (.I0(\slvo[3][hconfig][3] [23]),
        .I1(\slvo[2][hconfig][3] [23]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][3] [23]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][3] [23]),
        .O(\syncrregs.r[hrdatas][23]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][23]_i_25 
       (.I0(\slvo[7][hconfig][3] [23]),
        .I1(\slvo[6][hconfig][3] [23]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][3] [23]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][3] [23]),
        .O(\syncrregs.r[hrdatas][23]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][23]_i_26 
       (.I0(\slvo[3][hconfig][0] [23]),
        .I1(\slvo[2][hconfig][0] [23]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][0] [23]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][0] [23]),
        .O(\syncrregs.r[hrdatas][23]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][23]_i_27 
       (.I0(\slvo[7][hconfig][0] [23]),
        .I1(\slvo[6][hconfig][0] [23]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][0] [23]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][0] [23]),
        .O(\syncrregs.r[hrdatas][23]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][23]_i_28 
       (.I0(\slvo[3][hconfig][1] [23]),
        .I1(\slvo[2][hconfig][1] [23]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][1] [23]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][1] [23]),
        .O(\syncrregs.r[hrdatas][23]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][23]_i_29 
       (.I0(\slvo[7][hconfig][1] [23]),
        .I1(\slvo[6][hconfig][1] [23]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][1] [23]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][1] [23]),
        .O(\syncrregs.r[hrdatas][23]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][24]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][24]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][24]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][24]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][24]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][24]_i_14 
       (.I0(\slvo[3][hconfig][6] [24]),
        .I1(\slvo[2][hconfig][6] [24]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][6] [24]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][6] [24]),
        .O(\syncrregs.r[hrdatas][24]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][24]_i_15 
       (.I0(\slvo[7][hconfig][6] [24]),
        .I1(\slvo[6][hconfig][6] [24]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][6] [24]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][6] [24]),
        .O(\syncrregs.r[hrdatas][24]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][24]_i_16 
       (.I0(\slvo[3][hconfig][7] [24]),
        .I1(\slvo[2][hconfig][7] [24]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][7] [24]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][7] [24]),
        .O(\syncrregs.r[hrdatas][24]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][24]_i_17 
       (.I0(\slvo[7][hconfig][7] [24]),
        .I1(\slvo[6][hconfig][7] [24]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][7] [24]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][7] [24]),
        .O(\syncrregs.r[hrdatas][24]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][24]_i_18 
       (.I0(\slvo[3][hconfig][4] [24]),
        .I1(\slvo[2][hconfig][4] [24]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][4] [24]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][4] [24]),
        .O(\syncrregs.r[hrdatas][24]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][24]_i_19 
       (.I0(\slvo[7][hconfig][4] [24]),
        .I1(\slvo[6][hconfig][4] [24]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][4] [24]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][4] [24]),
        .O(\syncrregs.r[hrdatas][24]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][24]_i_20 
       (.I0(\slvo[3][hconfig][5] [24]),
        .I1(\slvo[2][hconfig][5] [24]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][5] [24]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][5] [24]),
        .O(\syncrregs.r[hrdatas][24]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][24]_i_21 
       (.I0(\slvo[7][hconfig][5] [24]),
        .I1(\slvo[6][hconfig][5] [24]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][5] [24]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][5] [24]),
        .O(\syncrregs.r[hrdatas][24]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][24]_i_22 
       (.I0(\slvo[3][hconfig][2] [24]),
        .I1(\slvo[2][hconfig][2] [24]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][2] [24]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][2] [24]),
        .O(\syncrregs.r[hrdatas][24]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][24]_i_23 
       (.I0(\slvo[7][hconfig][2] [24]),
        .I1(\slvo[6][hconfig][2] [24]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][2] [24]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][2] [24]),
        .O(\syncrregs.r[hrdatas][24]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][24]_i_24 
       (.I0(\slvo[3][hconfig][3] [24]),
        .I1(\slvo[2][hconfig][3] [24]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][3] [24]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][3] [24]),
        .O(\syncrregs.r[hrdatas][24]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][24]_i_25 
       (.I0(\slvo[7][hconfig][3] [24]),
        .I1(\slvo[6][hconfig][3] [24]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][3] [24]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][3] [24]),
        .O(\syncrregs.r[hrdatas][24]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][24]_i_26 
       (.I0(\slvo[3][hconfig][0] [24]),
        .I1(\slvo[2][hconfig][0] [24]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][0] [24]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][0] [24]),
        .O(\syncrregs.r[hrdatas][24]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][24]_i_27 
       (.I0(\slvo[7][hconfig][0] [24]),
        .I1(\slvo[6][hconfig][0] [24]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][0] [24]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][0] [24]),
        .O(\syncrregs.r[hrdatas][24]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][24]_i_28 
       (.I0(\slvo[3][hconfig][1] [24]),
        .I1(\slvo[2][hconfig][1] [24]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[1][hconfig][1] [24]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[0][hconfig][1] [24]),
        .O(\syncrregs.r[hrdatas][24]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][24]_i_29 
       (.I0(\slvo[7][hconfig][1] [24]),
        .I1(\slvo[6][hconfig][1] [24]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .I3(\slvo[5][hconfig][1] [24]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .I5(\slvo[4][hconfig][1] [24]),
        .O(\syncrregs.r[hrdatas][24]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][25]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][25]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][25]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][25]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][25]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][25]_i_14 
       (.I0(\slvo[3][hconfig][6] [25]),
        .I1(\slvo[2][hconfig][6] [25]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][6] [25]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][6] [25]),
        .O(\syncrregs.r[hrdatas][25]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][25]_i_15 
       (.I0(\slvo[7][hconfig][6] [25]),
        .I1(\slvo[6][hconfig][6] [25]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][6] [25]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][6] [25]),
        .O(\syncrregs.r[hrdatas][25]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][25]_i_16 
       (.I0(\slvo[3][hconfig][7] [25]),
        .I1(\slvo[2][hconfig][7] [25]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][7] [25]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][7] [25]),
        .O(\syncrregs.r[hrdatas][25]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][25]_i_17 
       (.I0(\slvo[7][hconfig][7] [25]),
        .I1(\slvo[6][hconfig][7] [25]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][7] [25]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][7] [25]),
        .O(\syncrregs.r[hrdatas][25]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][25]_i_18 
       (.I0(\slvo[3][hconfig][4] [25]),
        .I1(\slvo[2][hconfig][4] [25]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][4] [25]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][4] [25]),
        .O(\syncrregs.r[hrdatas][25]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][25]_i_19 
       (.I0(\slvo[7][hconfig][4] [25]),
        .I1(\slvo[6][hconfig][4] [25]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][4] [25]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][4] [25]),
        .O(\syncrregs.r[hrdatas][25]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][25]_i_20 
       (.I0(\slvo[3][hconfig][5] [25]),
        .I1(\slvo[2][hconfig][5] [25]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][5] [25]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][5] [25]),
        .O(\syncrregs.r[hrdatas][25]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][25]_i_21 
       (.I0(\slvo[7][hconfig][5] [25]),
        .I1(\slvo[6][hconfig][5] [25]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][5] [25]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][5] [25]),
        .O(\syncrregs.r[hrdatas][25]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][25]_i_22 
       (.I0(\slvo[3][hconfig][2] [25]),
        .I1(\slvo[2][hconfig][2] [25]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][2] [25]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][2] [25]),
        .O(\syncrregs.r[hrdatas][25]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][25]_i_23 
       (.I0(\slvo[7][hconfig][2] [25]),
        .I1(\slvo[6][hconfig][2] [25]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][2] [25]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][2] [25]),
        .O(\syncrregs.r[hrdatas][25]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][25]_i_24 
       (.I0(\slvo[3][hconfig][3] [25]),
        .I1(\slvo[2][hconfig][3] [25]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][3] [25]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][3] [25]),
        .O(\syncrregs.r[hrdatas][25]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][25]_i_25 
       (.I0(\slvo[7][hconfig][3] [25]),
        .I1(\slvo[6][hconfig][3] [25]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][3] [25]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][3] [25]),
        .O(\syncrregs.r[hrdatas][25]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][25]_i_26 
       (.I0(\slvo[3][hconfig][0] [25]),
        .I1(\slvo[2][hconfig][0] [25]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][0] [25]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][0] [25]),
        .O(\syncrregs.r[hrdatas][25]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][25]_i_27 
       (.I0(\slvo[7][hconfig][0] [25]),
        .I1(\slvo[6][hconfig][0] [25]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][0] [25]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][0] [25]),
        .O(\syncrregs.r[hrdatas][25]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][25]_i_28 
       (.I0(\slvo[3][hconfig][1] [25]),
        .I1(\slvo[2][hconfig][1] [25]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][1] [25]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][1] [25]),
        .O(\syncrregs.r[hrdatas][25]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][25]_i_29 
       (.I0(\slvo[7][hconfig][1] [25]),
        .I1(\slvo[6][hconfig][1] [25]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][1] [25]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][1] [25]),
        .O(\syncrregs.r[hrdatas][25]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][26]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][26]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][26]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][26]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][26]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][26]_i_14 
       (.I0(\slvo[3][hconfig][6] [26]),
        .I1(\slvo[2][hconfig][6] [26]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][6] [26]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][6] [26]),
        .O(\syncrregs.r[hrdatas][26]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][26]_i_15 
       (.I0(\slvo[7][hconfig][6] [26]),
        .I1(\slvo[6][hconfig][6] [26]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][6] [26]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][6] [26]),
        .O(\syncrregs.r[hrdatas][26]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][26]_i_16 
       (.I0(\slvo[3][hconfig][7] [26]),
        .I1(\slvo[2][hconfig][7] [26]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][7] [26]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][7] [26]),
        .O(\syncrregs.r[hrdatas][26]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][26]_i_17 
       (.I0(\slvo[7][hconfig][7] [26]),
        .I1(\slvo[6][hconfig][7] [26]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][7] [26]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][7] [26]),
        .O(\syncrregs.r[hrdatas][26]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][26]_i_18 
       (.I0(\slvo[3][hconfig][4] [26]),
        .I1(\slvo[2][hconfig][4] [26]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][4] [26]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][4] [26]),
        .O(\syncrregs.r[hrdatas][26]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][26]_i_19 
       (.I0(\slvo[7][hconfig][4] [26]),
        .I1(\slvo[6][hconfig][4] [26]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][4] [26]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][4] [26]),
        .O(\syncrregs.r[hrdatas][26]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][26]_i_20 
       (.I0(\slvo[3][hconfig][5] [26]),
        .I1(\slvo[2][hconfig][5] [26]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][5] [26]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][5] [26]),
        .O(\syncrregs.r[hrdatas][26]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][26]_i_21 
       (.I0(\slvo[7][hconfig][5] [26]),
        .I1(\slvo[6][hconfig][5] [26]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][5] [26]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][5] [26]),
        .O(\syncrregs.r[hrdatas][26]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][26]_i_22 
       (.I0(\slvo[3][hconfig][2] [26]),
        .I1(\slvo[2][hconfig][2] [26]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][2] [26]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][2] [26]),
        .O(\syncrregs.r[hrdatas][26]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][26]_i_23 
       (.I0(\slvo[7][hconfig][2] [26]),
        .I1(\slvo[6][hconfig][2] [26]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][2] [26]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][2] [26]),
        .O(\syncrregs.r[hrdatas][26]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][26]_i_24 
       (.I0(\slvo[3][hconfig][3] [26]),
        .I1(\slvo[2][hconfig][3] [26]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][3] [26]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][3] [26]),
        .O(\syncrregs.r[hrdatas][26]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][26]_i_25 
       (.I0(\slvo[7][hconfig][3] [26]),
        .I1(\slvo[6][hconfig][3] [26]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][3] [26]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][3] [26]),
        .O(\syncrregs.r[hrdatas][26]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][26]_i_26 
       (.I0(\slvo[3][hconfig][0] [26]),
        .I1(\slvo[2][hconfig][0] [26]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][0] [26]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][0] [26]),
        .O(\syncrregs.r[hrdatas][26]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][26]_i_27 
       (.I0(\slvo[7][hconfig][0] [26]),
        .I1(\slvo[6][hconfig][0] [26]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][0] [26]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][0] [26]),
        .O(\syncrregs.r[hrdatas][26]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][26]_i_28 
       (.I0(\slvo[3][hconfig][1] [26]),
        .I1(\slvo[2][hconfig][1] [26]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][1] [26]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][1] [26]),
        .O(\syncrregs.r[hrdatas][26]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][26]_i_29 
       (.I0(\slvo[7][hconfig][1] [26]),
        .I1(\slvo[6][hconfig][1] [26]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][1] [26]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][1] [26]),
        .O(\syncrregs.r[hrdatas][26]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][27]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][27]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][27]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][27]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][27]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][27]_i_14 
       (.I0(\slvo[3][hconfig][6] [27]),
        .I1(\slvo[2][hconfig][6] [27]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][6] [27]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][6] [27]),
        .O(\syncrregs.r[hrdatas][27]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][27]_i_15 
       (.I0(\slvo[7][hconfig][6] [27]),
        .I1(\slvo[6][hconfig][6] [27]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][6] [27]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][6] [27]),
        .O(\syncrregs.r[hrdatas][27]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][27]_i_16 
       (.I0(\slvo[3][hconfig][7] [27]),
        .I1(\slvo[2][hconfig][7] [27]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][7] [27]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][7] [27]),
        .O(\syncrregs.r[hrdatas][27]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][27]_i_17 
       (.I0(\slvo[7][hconfig][7] [27]),
        .I1(\slvo[6][hconfig][7] [27]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][7] [27]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][7] [27]),
        .O(\syncrregs.r[hrdatas][27]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][27]_i_18 
       (.I0(\slvo[3][hconfig][4] [27]),
        .I1(\slvo[2][hconfig][4] [27]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][4] [27]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][4] [27]),
        .O(\syncrregs.r[hrdatas][27]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][27]_i_19 
       (.I0(\slvo[7][hconfig][4] [27]),
        .I1(\slvo[6][hconfig][4] [27]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][4] [27]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][4] [27]),
        .O(\syncrregs.r[hrdatas][27]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][27]_i_20 
       (.I0(\slvo[3][hconfig][5] [27]),
        .I1(\slvo[2][hconfig][5] [27]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][5] [27]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][5] [27]),
        .O(\syncrregs.r[hrdatas][27]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][27]_i_21 
       (.I0(\slvo[7][hconfig][5] [27]),
        .I1(\slvo[6][hconfig][5] [27]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][5] [27]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][5] [27]),
        .O(\syncrregs.r[hrdatas][27]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][27]_i_22 
       (.I0(\slvo[3][hconfig][2] [27]),
        .I1(\slvo[2][hconfig][2] [27]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][2] [27]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][2] [27]),
        .O(\syncrregs.r[hrdatas][27]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][27]_i_23 
       (.I0(\slvo[7][hconfig][2] [27]),
        .I1(\slvo[6][hconfig][2] [27]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][2] [27]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][2] [27]),
        .O(\syncrregs.r[hrdatas][27]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][27]_i_24 
       (.I0(\slvo[3][hconfig][3] [27]),
        .I1(\slvo[2][hconfig][3] [27]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][3] [27]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][3] [27]),
        .O(\syncrregs.r[hrdatas][27]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][27]_i_25 
       (.I0(\slvo[7][hconfig][3] [27]),
        .I1(\slvo[6][hconfig][3] [27]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][3] [27]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][3] [27]),
        .O(\syncrregs.r[hrdatas][27]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][27]_i_26 
       (.I0(\slvo[3][hconfig][0] [27]),
        .I1(\slvo[2][hconfig][0] [27]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][0] [27]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][0] [27]),
        .O(\syncrregs.r[hrdatas][27]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][27]_i_27 
       (.I0(\slvo[7][hconfig][0] [27]),
        .I1(\slvo[6][hconfig][0] [27]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][0] [27]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][0] [27]),
        .O(\syncrregs.r[hrdatas][27]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][27]_i_28 
       (.I0(\slvo[3][hconfig][1] [27]),
        .I1(\slvo[2][hconfig][1] [27]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][1] [27]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][1] [27]),
        .O(\syncrregs.r[hrdatas][27]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][27]_i_29 
       (.I0(\slvo[7][hconfig][1] [27]),
        .I1(\slvo[6][hconfig][1] [27]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][1] [27]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][1] [27]),
        .O(\syncrregs.r[hrdatas][27]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][28]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][28]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][28]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][28]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][28]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][28]_i_14 
       (.I0(\slvo[3][hconfig][6] [28]),
        .I1(\slvo[2][hconfig][6] [28]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][6] [28]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][6] [28]),
        .O(\syncrregs.r[hrdatas][28]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][28]_i_15 
       (.I0(\slvo[7][hconfig][6] [28]),
        .I1(\slvo[6][hconfig][6] [28]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][6] [28]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][6] [28]),
        .O(\syncrregs.r[hrdatas][28]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][28]_i_16 
       (.I0(\slvo[3][hconfig][7] [28]),
        .I1(\slvo[2][hconfig][7] [28]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][7] [28]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][7] [28]),
        .O(\syncrregs.r[hrdatas][28]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][28]_i_17 
       (.I0(\slvo[7][hconfig][7] [28]),
        .I1(\slvo[6][hconfig][7] [28]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][7] [28]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][7] [28]),
        .O(\syncrregs.r[hrdatas][28]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][28]_i_18 
       (.I0(\slvo[3][hconfig][4] [28]),
        .I1(\slvo[2][hconfig][4] [28]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][4] [28]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][4] [28]),
        .O(\syncrregs.r[hrdatas][28]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][28]_i_19 
       (.I0(\slvo[7][hconfig][4] [28]),
        .I1(\slvo[6][hconfig][4] [28]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][4] [28]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][4] [28]),
        .O(\syncrregs.r[hrdatas][28]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][28]_i_20 
       (.I0(\slvo[3][hconfig][5] [28]),
        .I1(\slvo[2][hconfig][5] [28]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][5] [28]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][5] [28]),
        .O(\syncrregs.r[hrdatas][28]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][28]_i_21 
       (.I0(\slvo[7][hconfig][5] [28]),
        .I1(\slvo[6][hconfig][5] [28]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][5] [28]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][5] [28]),
        .O(\syncrregs.r[hrdatas][28]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][28]_i_22 
       (.I0(\slvo[3][hconfig][2] [28]),
        .I1(\slvo[2][hconfig][2] [28]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][2] [28]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][2] [28]),
        .O(\syncrregs.r[hrdatas][28]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][28]_i_23 
       (.I0(\slvo[7][hconfig][2] [28]),
        .I1(\slvo[6][hconfig][2] [28]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][2] [28]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][2] [28]),
        .O(\syncrregs.r[hrdatas][28]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][28]_i_24 
       (.I0(\slvo[3][hconfig][3] [28]),
        .I1(\slvo[2][hconfig][3] [28]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][3] [28]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][3] [28]),
        .O(\syncrregs.r[hrdatas][28]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][28]_i_25 
       (.I0(\slvo[7][hconfig][3] [28]),
        .I1(\slvo[6][hconfig][3] [28]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][3] [28]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][3] [28]),
        .O(\syncrregs.r[hrdatas][28]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][28]_i_26 
       (.I0(\slvo[3][hconfig][0] [28]),
        .I1(\slvo[2][hconfig][0] [28]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][0] [28]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][0] [28]),
        .O(\syncrregs.r[hrdatas][28]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][28]_i_27 
       (.I0(\slvo[7][hconfig][0] [28]),
        .I1(\slvo[6][hconfig][0] [28]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][0] [28]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][0] [28]),
        .O(\syncrregs.r[hrdatas][28]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][28]_i_28 
       (.I0(\slvo[3][hconfig][1] [28]),
        .I1(\slvo[2][hconfig][1] [28]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][1] [28]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][1] [28]),
        .O(\syncrregs.r[hrdatas][28]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][28]_i_29 
       (.I0(\slvo[7][hconfig][1] [28]),
        .I1(\slvo[6][hconfig][1] [28]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][1] [28]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][1] [28]),
        .O(\syncrregs.r[hrdatas][28]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][29]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][29]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][29]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][29]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][29]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][29]_i_14 
       (.I0(\slvo[3][hconfig][6] [29]),
        .I1(\slvo[2][hconfig][6] [29]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][6] [29]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][6] [29]),
        .O(\syncrregs.r[hrdatas][29]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][29]_i_15 
       (.I0(\slvo[7][hconfig][6] [29]),
        .I1(\slvo[6][hconfig][6] [29]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][6] [29]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][6] [29]),
        .O(\syncrregs.r[hrdatas][29]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][29]_i_16 
       (.I0(\slvo[3][hconfig][7] [29]),
        .I1(\slvo[2][hconfig][7] [29]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][7] [29]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][7] [29]),
        .O(\syncrregs.r[hrdatas][29]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][29]_i_17 
       (.I0(\slvo[7][hconfig][7] [29]),
        .I1(\slvo[6][hconfig][7] [29]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][7] [29]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][7] [29]),
        .O(\syncrregs.r[hrdatas][29]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][29]_i_18 
       (.I0(\slvo[3][hconfig][4] [29]),
        .I1(\slvo[2][hconfig][4] [29]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][4] [29]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][4] [29]),
        .O(\syncrregs.r[hrdatas][29]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][29]_i_19 
       (.I0(\slvo[7][hconfig][4] [29]),
        .I1(\slvo[6][hconfig][4] [29]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][4] [29]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][4] [29]),
        .O(\syncrregs.r[hrdatas][29]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][29]_i_20 
       (.I0(\slvo[3][hconfig][5] [29]),
        .I1(\slvo[2][hconfig][5] [29]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][5] [29]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][5] [29]),
        .O(\syncrregs.r[hrdatas][29]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][29]_i_21 
       (.I0(\slvo[7][hconfig][5] [29]),
        .I1(\slvo[6][hconfig][5] [29]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][5] [29]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][5] [29]),
        .O(\syncrregs.r[hrdatas][29]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][29]_i_22 
       (.I0(\slvo[3][hconfig][2] [29]),
        .I1(\slvo[2][hconfig][2] [29]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][2] [29]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][2] [29]),
        .O(\syncrregs.r[hrdatas][29]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][29]_i_23 
       (.I0(\slvo[7][hconfig][2] [29]),
        .I1(\slvo[6][hconfig][2] [29]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][2] [29]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][2] [29]),
        .O(\syncrregs.r[hrdatas][29]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][29]_i_24 
       (.I0(\slvo[3][hconfig][3] [29]),
        .I1(\slvo[2][hconfig][3] [29]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][3] [29]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][3] [29]),
        .O(\syncrregs.r[hrdatas][29]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][29]_i_25 
       (.I0(\slvo[7][hconfig][3] [29]),
        .I1(\slvo[6][hconfig][3] [29]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][3] [29]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][3] [29]),
        .O(\syncrregs.r[hrdatas][29]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][29]_i_26 
       (.I0(\slvo[3][hconfig][0] [29]),
        .I1(\slvo[2][hconfig][0] [29]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][0] [29]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][0] [29]),
        .O(\syncrregs.r[hrdatas][29]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][29]_i_27 
       (.I0(\slvo[7][hconfig][0] [29]),
        .I1(\slvo[6][hconfig][0] [29]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][0] [29]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][0] [29]),
        .O(\syncrregs.r[hrdatas][29]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][29]_i_28 
       (.I0(\slvo[3][hconfig][1] [29]),
        .I1(\slvo[2][hconfig][1] [29]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][1] [29]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][1] [29]),
        .O(\syncrregs.r[hrdatas][29]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][29]_i_29 
       (.I0(\slvo[7][hconfig][1] [29]),
        .I1(\slvo[6][hconfig][1] [29]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][1] [29]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][1] [29]),
        .O(\syncrregs.r[hrdatas][29]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][2]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][2]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][2]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][2]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][2]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][2]_i_14 
       (.I0(\slvo[3][hconfig][6] [2]),
        .I1(\slvo[2][hconfig][6] [2]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][6] [2]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][6] [2]),
        .O(\syncrregs.r[hrdatas][2]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][2]_i_15 
       (.I0(\slvo[7][hconfig][6] [2]),
        .I1(\slvo[6][hconfig][6] [2]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][6] [2]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][6] [2]),
        .O(\syncrregs.r[hrdatas][2]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][2]_i_16 
       (.I0(\slvo[3][hconfig][7] [2]),
        .I1(\slvo[2][hconfig][7] [2]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][7] [2]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][7] [2]),
        .O(\syncrregs.r[hrdatas][2]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][2]_i_17 
       (.I0(\slvo[7][hconfig][7] [2]),
        .I1(\slvo[6][hconfig][7] [2]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][7] [2]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][7] [2]),
        .O(\syncrregs.r[hrdatas][2]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][2]_i_18 
       (.I0(\slvo[3][hconfig][4] [2]),
        .I1(\slvo[2][hconfig][4] [2]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][4] [2]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][4] [2]),
        .O(\syncrregs.r[hrdatas][2]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][2]_i_19 
       (.I0(\slvo[7][hconfig][4] [2]),
        .I1(\slvo[6][hconfig][4] [2]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][4] [2]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][4] [2]),
        .O(\syncrregs.r[hrdatas][2]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][2]_i_20 
       (.I0(\slvo[3][hconfig][5] [2]),
        .I1(\slvo[2][hconfig][5] [2]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][5] [2]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][5] [2]),
        .O(\syncrregs.r[hrdatas][2]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][2]_i_21 
       (.I0(\slvo[7][hconfig][5] [2]),
        .I1(\slvo[6][hconfig][5] [2]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][5] [2]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][5] [2]),
        .O(\syncrregs.r[hrdatas][2]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][2]_i_22 
       (.I0(\slvo[3][hconfig][2] [2]),
        .I1(\slvo[2][hconfig][2] [2]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][2] [2]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][2] [2]),
        .O(\syncrregs.r[hrdatas][2]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][2]_i_23 
       (.I0(\slvo[7][hconfig][2] [2]),
        .I1(\slvo[6][hconfig][2] [2]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][2] [2]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][2] [2]),
        .O(\syncrregs.r[hrdatas][2]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][2]_i_24 
       (.I0(\slvo[3][hconfig][3] [2]),
        .I1(\slvo[2][hconfig][3] [2]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][3] [2]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][3] [2]),
        .O(\syncrregs.r[hrdatas][2]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][2]_i_25 
       (.I0(\slvo[7][hconfig][3] [2]),
        .I1(\slvo[6][hconfig][3] [2]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][3] [2]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][3] [2]),
        .O(\syncrregs.r[hrdatas][2]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][2]_i_26 
       (.I0(\slvo[3][hconfig][0] [2]),
        .I1(\slvo[2][hconfig][0] [2]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][0] [2]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][0] [2]),
        .O(\syncrregs.r[hrdatas][2]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][2]_i_27 
       (.I0(\slvo[7][hconfig][0] [2]),
        .I1(\slvo[6][hconfig][0] [2]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][0] [2]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][0] [2]),
        .O(\syncrregs.r[hrdatas][2]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][2]_i_28 
       (.I0(\slvo[3][hconfig][1] [2]),
        .I1(\slvo[2][hconfig][1] [2]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][1] [2]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][1] [2]),
        .O(\syncrregs.r[hrdatas][2]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][2]_i_29 
       (.I0(\slvo[7][hconfig][1] [2]),
        .I1(\slvo[6][hconfig][1] [2]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][1] [2]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][1] [2]),
        .O(\syncrregs.r[hrdatas][2]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][30]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][30]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][30]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][30]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][30]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][30]_i_14 
       (.I0(\slvo[3][hconfig][6] [30]),
        .I1(\slvo[2][hconfig][6] [30]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][6] [30]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][6] [30]),
        .O(\syncrregs.r[hrdatas][30]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][30]_i_15 
       (.I0(\slvo[7][hconfig][6] [30]),
        .I1(\slvo[6][hconfig][6] [30]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][6] [30]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][6] [30]),
        .O(\syncrregs.r[hrdatas][30]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][30]_i_16 
       (.I0(\slvo[3][hconfig][7] [30]),
        .I1(\slvo[2][hconfig][7] [30]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][7] [30]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][7] [30]),
        .O(\syncrregs.r[hrdatas][30]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][30]_i_17 
       (.I0(\slvo[7][hconfig][7] [30]),
        .I1(\slvo[6][hconfig][7] [30]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][7] [30]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][7] [30]),
        .O(\syncrregs.r[hrdatas][30]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][30]_i_18 
       (.I0(\slvo[3][hconfig][4] [30]),
        .I1(\slvo[2][hconfig][4] [30]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][4] [30]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][4] [30]),
        .O(\syncrregs.r[hrdatas][30]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][30]_i_19 
       (.I0(\slvo[7][hconfig][4] [30]),
        .I1(\slvo[6][hconfig][4] [30]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][4] [30]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][4] [30]),
        .O(\syncrregs.r[hrdatas][30]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][30]_i_20 
       (.I0(\slvo[3][hconfig][5] [30]),
        .I1(\slvo[2][hconfig][5] [30]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][5] [30]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][5] [30]),
        .O(\syncrregs.r[hrdatas][30]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][30]_i_21 
       (.I0(\slvo[7][hconfig][5] [30]),
        .I1(\slvo[6][hconfig][5] [30]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][5] [30]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][5] [30]),
        .O(\syncrregs.r[hrdatas][30]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][30]_i_22 
       (.I0(\slvo[3][hconfig][2] [30]),
        .I1(\slvo[2][hconfig][2] [30]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][2] [30]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][2] [30]),
        .O(\syncrregs.r[hrdatas][30]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][30]_i_23 
       (.I0(\slvo[7][hconfig][2] [30]),
        .I1(\slvo[6][hconfig][2] [30]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][2] [30]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][2] [30]),
        .O(\syncrregs.r[hrdatas][30]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][30]_i_24 
       (.I0(\slvo[3][hconfig][3] [30]),
        .I1(\slvo[2][hconfig][3] [30]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][3] [30]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][3] [30]),
        .O(\syncrregs.r[hrdatas][30]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][30]_i_25 
       (.I0(\slvo[7][hconfig][3] [30]),
        .I1(\slvo[6][hconfig][3] [30]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][3] [30]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][3] [30]),
        .O(\syncrregs.r[hrdatas][30]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][30]_i_26 
       (.I0(\slvo[3][hconfig][0] [30]),
        .I1(\slvo[2][hconfig][0] [30]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][0] [30]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][0] [30]),
        .O(\syncrregs.r[hrdatas][30]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][30]_i_27 
       (.I0(\slvo[7][hconfig][0] [30]),
        .I1(\slvo[6][hconfig][0] [30]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][0] [30]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][0] [30]),
        .O(\syncrregs.r[hrdatas][30]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][30]_i_28 
       (.I0(\slvo[3][hconfig][1] [30]),
        .I1(\slvo[2][hconfig][1] [30]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][1] [30]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][1] [30]),
        .O(\syncrregs.r[hrdatas][30]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][30]_i_29 
       (.I0(\slvo[7][hconfig][1] [30]),
        .I1(\slvo[6][hconfig][1] [30]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][1] [30]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][1] [30]),
        .O(\syncrregs.r[hrdatas][30]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h80000000F7FFFFFF)) 
    \syncrregs.r[hrdatas][31]_i_1 
       (.I0(sel0[4]),
        .I1(sel0[5]),
        .I2(\syncrregs.r[hrdatas][31]_i_3_n_0 ),
        .I3(sel0[3]),
        .I4(sel0[6]),
        .I5(p_179_out),
        .O(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][31]_i_17 
       (.I0(\slvo[3][hconfig][6] [31]),
        .I1(\slvo[2][hconfig][6] [31]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][6] [31]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][6] [31]),
        .O(\syncrregs.r[hrdatas][31]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][31]_i_18 
       (.I0(\slvo[7][hconfig][6] [31]),
        .I1(\slvo[6][hconfig][6] [31]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][6] [31]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][6] [31]),
        .O(\syncrregs.r[hrdatas][31]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][31]_i_19 
       (.I0(\slvo[3][hconfig][7] [31]),
        .I1(\slvo[2][hconfig][7] [31]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][7] [31]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][7] [31]),
        .O(\syncrregs.r[hrdatas][31]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][31]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][31]_i_5_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][31]_i_6_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][31]_i_7_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][31]_i_8_n_0 ),
        .O(\slvo[15][hready]__0 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][31]_i_20 
       (.I0(\slvo[7][hconfig][7] [31]),
        .I1(\slvo[6][hconfig][7] [31]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][7] [31]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][7] [31]),
        .O(\syncrregs.r[hrdatas][31]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][31]_i_21 
       (.I0(\slvo[3][hconfig][4] [31]),
        .I1(\slvo[2][hconfig][4] [31]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][4] [31]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][4] [31]),
        .O(\syncrregs.r[hrdatas][31]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][31]_i_22 
       (.I0(\slvo[7][hconfig][4] [31]),
        .I1(\slvo[6][hconfig][4] [31]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][4] [31]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][4] [31]),
        .O(\syncrregs.r[hrdatas][31]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][31]_i_23 
       (.I0(\slvo[3][hconfig][5] [31]),
        .I1(\slvo[2][hconfig][5] [31]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][5] [31]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][5] [31]),
        .O(\syncrregs.r[hrdatas][31]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][31]_i_24 
       (.I0(\slvo[7][hconfig][5] [31]),
        .I1(\slvo[6][hconfig][5] [31]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][5] [31]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][5] [31]),
        .O(\syncrregs.r[hrdatas][31]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][31]_i_25 
       (.I0(\slvo[3][hconfig][2] [31]),
        .I1(\slvo[2][hconfig][2] [31]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][2] [31]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][2] [31]),
        .O(\syncrregs.r[hrdatas][31]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][31]_i_26 
       (.I0(\slvo[7][hconfig][2] [31]),
        .I1(\slvo[6][hconfig][2] [31]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][2] [31]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][2] [31]),
        .O(\syncrregs.r[hrdatas][31]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][31]_i_27 
       (.I0(\slvo[3][hconfig][3] [31]),
        .I1(\slvo[2][hconfig][3] [31]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][3] [31]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][3] [31]),
        .O(\syncrregs.r[hrdatas][31]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][31]_i_28 
       (.I0(\slvo[7][hconfig][3] [31]),
        .I1(\slvo[6][hconfig][3] [31]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][3] [31]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][3] [31]),
        .O(\syncrregs.r[hrdatas][31]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][31]_i_29 
       (.I0(\slvo[3][hconfig][0] [31]),
        .I1(\slvo[2][hconfig][0] [31]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][0] [31]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][0] [31]),
        .O(\syncrregs.r[hrdatas][31]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h80FF)) 
    \syncrregs.r[hrdatas][31]_i_3 
       (.I0(sel0[1]),
        .I1(sel0[2]),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(p_179_out),
        .O(\syncrregs.r[hrdatas][31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][31]_i_30 
       (.I0(\slvo[7][hconfig][0] [31]),
        .I1(\slvo[6][hconfig][0] [31]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][0] [31]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][0] [31]),
        .O(\syncrregs.r[hrdatas][31]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][31]_i_31 
       (.I0(\slvo[3][hconfig][1] [31]),
        .I1(\slvo[2][hconfig][1] [31]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[1][hconfig][1] [31]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[0][hconfig][1] [31]),
        .O(\syncrregs.r[hrdatas][31]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][31]_i_32 
       (.I0(\slvo[7][hconfig][1] [31]),
        .I1(\slvo[6][hconfig][1] [31]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .I3(\slvo[5][hconfig][1] [31]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .I5(\slvo[4][hconfig][1] [31]),
        .O(\syncrregs.r[hrdatas][31]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0100010001000101)) 
    \syncrregs.r[hrdatas][31]_i_4 
       (.I0(sel0[5]),
        .I1(sel0[4]),
        .I2(sel0[6]),
        .I3(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I4(\syncrregs.r_reg[haddr_n_0_][2] ),
        .I5(\syncrregs.r_reg[haddr_n_0_][3] ),
        .O(p_179_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][3]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][3]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][3]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][3]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][3]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][3]_i_14 
       (.I0(\slvo[3][hconfig][6] [3]),
        .I1(\slvo[2][hconfig][6] [3]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][6] [3]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][6] [3]),
        .O(\syncrregs.r[hrdatas][3]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][3]_i_15 
       (.I0(\slvo[7][hconfig][6] [3]),
        .I1(\slvo[6][hconfig][6] [3]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][6] [3]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][6] [3]),
        .O(\syncrregs.r[hrdatas][3]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][3]_i_16 
       (.I0(\slvo[3][hconfig][7] [3]),
        .I1(\slvo[2][hconfig][7] [3]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][7] [3]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][7] [3]),
        .O(\syncrregs.r[hrdatas][3]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][3]_i_17 
       (.I0(\slvo[7][hconfig][7] [3]),
        .I1(\slvo[6][hconfig][7] [3]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][7] [3]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][7] [3]),
        .O(\syncrregs.r[hrdatas][3]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][3]_i_18 
       (.I0(\slvo[3][hconfig][4] [3]),
        .I1(\slvo[2][hconfig][4] [3]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][4] [3]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][4] [3]),
        .O(\syncrregs.r[hrdatas][3]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][3]_i_19 
       (.I0(\slvo[7][hconfig][4] [3]),
        .I1(\slvo[6][hconfig][4] [3]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][4] [3]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][4] [3]),
        .O(\syncrregs.r[hrdatas][3]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][3]_i_20 
       (.I0(\slvo[3][hconfig][5] [3]),
        .I1(\slvo[2][hconfig][5] [3]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][5] [3]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][5] [3]),
        .O(\syncrregs.r[hrdatas][3]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][3]_i_21 
       (.I0(\slvo[7][hconfig][5] [3]),
        .I1(\slvo[6][hconfig][5] [3]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][5] [3]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][5] [3]),
        .O(\syncrregs.r[hrdatas][3]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][3]_i_22 
       (.I0(\slvo[3][hconfig][2] [3]),
        .I1(\slvo[2][hconfig][2] [3]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][2] [3]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][2] [3]),
        .O(\syncrregs.r[hrdatas][3]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][3]_i_23 
       (.I0(\slvo[7][hconfig][2] [3]),
        .I1(\slvo[6][hconfig][2] [3]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][2] [3]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][2] [3]),
        .O(\syncrregs.r[hrdatas][3]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][3]_i_24 
       (.I0(\slvo[3][hconfig][3] [3]),
        .I1(\slvo[2][hconfig][3] [3]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][3] [3]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][3] [3]),
        .O(\syncrregs.r[hrdatas][3]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][3]_i_25 
       (.I0(\slvo[7][hconfig][3] [3]),
        .I1(\slvo[6][hconfig][3] [3]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][3] [3]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][3] [3]),
        .O(\syncrregs.r[hrdatas][3]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][3]_i_26 
       (.I0(\slvo[3][hconfig][0] [3]),
        .I1(\slvo[2][hconfig][0] [3]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][0] [3]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][0] [3]),
        .O(\syncrregs.r[hrdatas][3]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][3]_i_27 
       (.I0(\slvo[7][hconfig][0] [3]),
        .I1(\slvo[6][hconfig][0] [3]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][0] [3]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][0] [3]),
        .O(\syncrregs.r[hrdatas][3]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][3]_i_28 
       (.I0(\slvo[3][hconfig][1] [3]),
        .I1(\slvo[2][hconfig][1] [3]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][1] [3]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][1] [3]),
        .O(\syncrregs.r[hrdatas][3]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][3]_i_29 
       (.I0(\slvo[7][hconfig][1] [3]),
        .I1(\slvo[6][hconfig][1] [3]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][1] [3]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][1] [3]),
        .O(\syncrregs.r[hrdatas][3]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][4]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][4]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][4]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][4]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][4]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][4]_i_14 
       (.I0(\slvo[3][hconfig][6] [4]),
        .I1(\slvo[2][hconfig][6] [4]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][6] [4]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][6] [4]),
        .O(\syncrregs.r[hrdatas][4]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][4]_i_15 
       (.I0(\slvo[7][hconfig][6] [4]),
        .I1(\slvo[6][hconfig][6] [4]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][6] [4]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][6] [4]),
        .O(\syncrregs.r[hrdatas][4]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][4]_i_16 
       (.I0(\slvo[3][hconfig][7] [4]),
        .I1(\slvo[2][hconfig][7] [4]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][7] [4]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][7] [4]),
        .O(\syncrregs.r[hrdatas][4]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][4]_i_17 
       (.I0(\slvo[7][hconfig][7] [4]),
        .I1(\slvo[6][hconfig][7] [4]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][7] [4]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][7] [4]),
        .O(\syncrregs.r[hrdatas][4]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][4]_i_18 
       (.I0(\slvo[3][hconfig][4] [4]),
        .I1(\slvo[2][hconfig][4] [4]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][4] [4]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][4] [4]),
        .O(\syncrregs.r[hrdatas][4]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][4]_i_19 
       (.I0(\slvo[7][hconfig][4] [4]),
        .I1(\slvo[6][hconfig][4] [4]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][4] [4]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][4] [4]),
        .O(\syncrregs.r[hrdatas][4]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][4]_i_20 
       (.I0(\slvo[3][hconfig][5] [4]),
        .I1(\slvo[2][hconfig][5] [4]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][5] [4]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][5] [4]),
        .O(\syncrregs.r[hrdatas][4]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][4]_i_21 
       (.I0(\slvo[7][hconfig][5] [4]),
        .I1(\slvo[6][hconfig][5] [4]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][5] [4]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][5] [4]),
        .O(\syncrregs.r[hrdatas][4]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][4]_i_22 
       (.I0(\slvo[3][hconfig][2] [4]),
        .I1(\slvo[2][hconfig][2] [4]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][2] [4]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][2] [4]),
        .O(\syncrregs.r[hrdatas][4]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][4]_i_23 
       (.I0(\slvo[7][hconfig][2] [4]),
        .I1(\slvo[6][hconfig][2] [4]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][2] [4]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][2] [4]),
        .O(\syncrregs.r[hrdatas][4]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][4]_i_24 
       (.I0(\slvo[3][hconfig][3] [4]),
        .I1(\slvo[2][hconfig][3] [4]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][3] [4]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][3] [4]),
        .O(\syncrregs.r[hrdatas][4]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][4]_i_25 
       (.I0(\slvo[7][hconfig][3] [4]),
        .I1(\slvo[6][hconfig][3] [4]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][3] [4]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][3] [4]),
        .O(\syncrregs.r[hrdatas][4]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][4]_i_26 
       (.I0(\slvo[3][hconfig][0] [4]),
        .I1(\slvo[2][hconfig][0] [4]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][0] [4]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][0] [4]),
        .O(\syncrregs.r[hrdatas][4]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][4]_i_27 
       (.I0(\slvo[7][hconfig][0] [4]),
        .I1(\slvo[6][hconfig][0] [4]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][0] [4]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][0] [4]),
        .O(\syncrregs.r[hrdatas][4]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][4]_i_28 
       (.I0(\slvo[3][hconfig][1] [4]),
        .I1(\slvo[2][hconfig][1] [4]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][1] [4]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][1] [4]),
        .O(\syncrregs.r[hrdatas][4]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][4]_i_29 
       (.I0(\slvo[7][hconfig][1] [4]),
        .I1(\slvo[6][hconfig][1] [4]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][1] [4]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][1] [4]),
        .O(\syncrregs.r[hrdatas][4]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEE222E200000000)) 
    \syncrregs.r[hrdatas][5]_i_1 
       (.I0(\syncrregs.r[hrdatas][5]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I2(\syncrregs.r_reg[hrdatas][5]_i_3_n_0 ),
        .I3(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I4(\syncrregs.r_reg[hrdatas][5]_i_4_n_0 ),
        .I5(p_179_out),
        .O(\syncrregs.r[hrdatas][5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][5]_i_13 
       (.I0(\slvo[3][hconfig][3] [5]),
        .I1(\slvo[2][hconfig][3] [5]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][3] [5]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][3] [5]),
        .O(\syncrregs.r[hrdatas][5]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][5]_i_14 
       (.I0(\slvo[7][hconfig][3] [5]),
        .I1(\slvo[6][hconfig][3] [5]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][3] [5]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][3] [5]),
        .O(\syncrregs.r[hrdatas][5]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][5]_i_15 
       (.I0(\slvo[3][hconfig][2] [5]),
        .I1(\slvo[2][hconfig][2] [5]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][2] [5]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][2] [5]),
        .O(\syncrregs.r[hrdatas][5]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][5]_i_16 
       (.I0(\slvo[7][hconfig][2] [5]),
        .I1(\slvo[6][hconfig][2] [5]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][2] [5]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][2] [5]),
        .O(\syncrregs.r[hrdatas][5]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][5]_i_17 
       (.I0(\slvo[3][hconfig][1] [5]),
        .I1(\slvo[2][hconfig][1] [5]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][1] [5]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][1] [5]),
        .O(\syncrregs.r[hrdatas][5]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][5]_i_18 
       (.I0(\slvo[7][hconfig][1] [5]),
        .I1(\slvo[6][hconfig][1] [5]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][1] [5]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][1] [5]),
        .O(\syncrregs.r[hrdatas][5]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][5]_i_19 
       (.I0(\slvo[3][hconfig][0] [5]),
        .I1(\slvo[2][hconfig][0] [5]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][0] [5]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][0] [5]),
        .O(\syncrregs.r[hrdatas][5]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][5]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][5]_i_5_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][5]_i_6_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I3(\syncrregs.r_reg[hrdatas][5]_i_7_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][2] ),
        .I5(\syncrregs.r_reg[hrdatas][5]_i_8_n_0 ),
        .O(\syncrregs.r[hrdatas][5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][5]_i_20 
       (.I0(\slvo[7][hconfig][0] [5]),
        .I1(\slvo[6][hconfig][0] [5]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][0] [5]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][0] [5]),
        .O(\syncrregs.r[hrdatas][5]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][5]_i_21 
       (.I0(\slvo[3][hconfig][4] [5]),
        .I1(\slvo[2][hconfig][4] [5]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][4] [5]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][4] [5]),
        .O(\syncrregs.r[hrdatas][5]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][5]_i_22 
       (.I0(\slvo[7][hconfig][4] [5]),
        .I1(\slvo[6][hconfig][4] [5]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][4] [5]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][4] [5]),
        .O(\syncrregs.r[hrdatas][5]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][5]_i_23 
       (.I0(\slvo[3][hconfig][5] [5]),
        .I1(\slvo[2][hconfig][5] [5]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][5] [5]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][5] [5]),
        .O(\syncrregs.r[hrdatas][5]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][5]_i_24 
       (.I0(\slvo[7][hconfig][5] [5]),
        .I1(\slvo[6][hconfig][5] [5]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][5] [5]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][5] [5]),
        .O(\syncrregs.r[hrdatas][5]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][5]_i_25 
       (.I0(\slvo[3][hconfig][6] [5]),
        .I1(\slvo[2][hconfig][6] [5]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][6] [5]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][6] [5]),
        .O(\syncrregs.r[hrdatas][5]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][5]_i_26 
       (.I0(\slvo[7][hconfig][6] [5]),
        .I1(\slvo[6][hconfig][6] [5]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][6] [5]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][6] [5]),
        .O(\syncrregs.r[hrdatas][5]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][5]_i_27 
       (.I0(\slvo[3][hconfig][7] [5]),
        .I1(\slvo[2][hconfig][7] [5]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][7] [5]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][7] [5]),
        .O(\syncrregs.r[hrdatas][5]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][5]_i_28 
       (.I0(\slvo[7][hconfig][7] [5]),
        .I1(\slvo[6][hconfig][7] [5]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][7] [5]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][7] [5]),
        .O(\syncrregs.r[hrdatas][5]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEE222E200000000)) 
    \syncrregs.r[hrdatas][6]_i_1 
       (.I0(\syncrregs.r[hrdatas][6]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I2(\syncrregs.r_reg[hrdatas][6]_i_3_n_0 ),
        .I3(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I4(\syncrregs.r_reg[hrdatas][6]_i_4_n_0 ),
        .I5(p_179_out),
        .O(\syncrregs.r[hrdatas][6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][6]_i_13 
       (.I0(\slvo[3][hconfig][3] [6]),
        .I1(\slvo[2][hconfig][3] [6]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][3] [6]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][3] [6]),
        .O(\syncrregs.r[hrdatas][6]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][6]_i_14 
       (.I0(\slvo[7][hconfig][3] [6]),
        .I1(\slvo[6][hconfig][3] [6]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][3] [6]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][3] [6]),
        .O(\syncrregs.r[hrdatas][6]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][6]_i_15 
       (.I0(\slvo[3][hconfig][2] [6]),
        .I1(\slvo[2][hconfig][2] [6]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][2] [6]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][2] [6]),
        .O(\syncrregs.r[hrdatas][6]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][6]_i_16 
       (.I0(\slvo[7][hconfig][2] [6]),
        .I1(\slvo[6][hconfig][2] [6]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][2] [6]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][2] [6]),
        .O(\syncrregs.r[hrdatas][6]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][6]_i_17 
       (.I0(\slvo[3][hconfig][1] [6]),
        .I1(\slvo[2][hconfig][1] [6]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][1] [6]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][1] [6]),
        .O(\syncrregs.r[hrdatas][6]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][6]_i_18 
       (.I0(\slvo[7][hconfig][1] [6]),
        .I1(\slvo[6][hconfig][1] [6]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][1] [6]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][1] [6]),
        .O(\syncrregs.r[hrdatas][6]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][6]_i_19 
       (.I0(\slvo[3][hconfig][0] [6]),
        .I1(\slvo[2][hconfig][0] [6]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][0] [6]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][0] [6]),
        .O(\syncrregs.r[hrdatas][6]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][6]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][6]_i_5_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][6]_i_6_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I3(\syncrregs.r_reg[hrdatas][6]_i_7_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][2] ),
        .I5(\syncrregs.r_reg[hrdatas][6]_i_8_n_0 ),
        .O(\syncrregs.r[hrdatas][6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][6]_i_20 
       (.I0(\slvo[7][hconfig][0] [6]),
        .I1(\slvo[6][hconfig][0] [6]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][0] [6]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][0] [6]),
        .O(\syncrregs.r[hrdatas][6]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][6]_i_21 
       (.I0(\slvo[3][hconfig][4] [6]),
        .I1(\slvo[2][hconfig][4] [6]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][4] [6]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][4] [6]),
        .O(\syncrregs.r[hrdatas][6]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][6]_i_22 
       (.I0(\slvo[7][hconfig][4] [6]),
        .I1(\slvo[6][hconfig][4] [6]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][4] [6]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][4] [6]),
        .O(\syncrregs.r[hrdatas][6]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][6]_i_23 
       (.I0(\slvo[3][hconfig][5] [6]),
        .I1(\slvo[2][hconfig][5] [6]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][5] [6]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][5] [6]),
        .O(\syncrregs.r[hrdatas][6]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][6]_i_24 
       (.I0(\slvo[7][hconfig][5] [6]),
        .I1(\slvo[6][hconfig][5] [6]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][5] [6]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][5] [6]),
        .O(\syncrregs.r[hrdatas][6]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][6]_i_25 
       (.I0(\slvo[3][hconfig][6] [6]),
        .I1(\slvo[2][hconfig][6] [6]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][6] [6]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][6] [6]),
        .O(\syncrregs.r[hrdatas][6]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][6]_i_26 
       (.I0(\slvo[7][hconfig][6] [6]),
        .I1(\slvo[6][hconfig][6] [6]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][6] [6]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][6] [6]),
        .O(\syncrregs.r[hrdatas][6]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][6]_i_27 
       (.I0(\slvo[3][hconfig][7] [6]),
        .I1(\slvo[2][hconfig][7] [6]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[1][hconfig][7] [6]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[0][hconfig][7] [6]),
        .O(\syncrregs.r[hrdatas][6]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][6]_i_28 
       (.I0(\slvo[7][hconfig][7] [6]),
        .I1(\slvo[6][hconfig][7] [6]),
        .I2(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .I3(\slvo[5][hconfig][7] [6]),
        .I4(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .I5(\slvo[4][hconfig][7] [6]),
        .O(\syncrregs.r[hrdatas][6]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][7]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][7]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][7]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][7]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][7]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][7]_i_14 
       (.I0(\slvo[3][hconfig][6] [7]),
        .I1(\slvo[2][hconfig][6] [7]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][6] [7]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][6] [7]),
        .O(\syncrregs.r[hrdatas][7]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][7]_i_15 
       (.I0(\slvo[7][hconfig][6] [7]),
        .I1(\slvo[6][hconfig][6] [7]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][6] [7]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][6] [7]),
        .O(\syncrregs.r[hrdatas][7]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][7]_i_16 
       (.I0(\slvo[3][hconfig][7] [7]),
        .I1(\slvo[2][hconfig][7] [7]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][7] [7]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][7] [7]),
        .O(\syncrregs.r[hrdatas][7]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][7]_i_17 
       (.I0(\slvo[7][hconfig][7] [7]),
        .I1(\slvo[6][hconfig][7] [7]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][7] [7]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][7] [7]),
        .O(\syncrregs.r[hrdatas][7]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][7]_i_18 
       (.I0(\slvo[3][hconfig][4] [7]),
        .I1(\slvo[2][hconfig][4] [7]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][4] [7]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][4] [7]),
        .O(\syncrregs.r[hrdatas][7]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][7]_i_19 
       (.I0(\slvo[7][hconfig][4] [7]),
        .I1(\slvo[6][hconfig][4] [7]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][4] [7]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][4] [7]),
        .O(\syncrregs.r[hrdatas][7]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][7]_i_20 
       (.I0(\slvo[3][hconfig][5] [7]),
        .I1(\slvo[2][hconfig][5] [7]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][5] [7]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][5] [7]),
        .O(\syncrregs.r[hrdatas][7]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][7]_i_21 
       (.I0(\slvo[7][hconfig][5] [7]),
        .I1(\slvo[6][hconfig][5] [7]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][5] [7]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][5] [7]),
        .O(\syncrregs.r[hrdatas][7]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][7]_i_22 
       (.I0(\slvo[3][hconfig][2] [7]),
        .I1(\slvo[2][hconfig][2] [7]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][2] [7]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][2] [7]),
        .O(\syncrregs.r[hrdatas][7]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][7]_i_23 
       (.I0(\slvo[7][hconfig][2] [7]),
        .I1(\slvo[6][hconfig][2] [7]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][2] [7]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][2] [7]),
        .O(\syncrregs.r[hrdatas][7]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][7]_i_24 
       (.I0(\slvo[3][hconfig][3] [7]),
        .I1(\slvo[2][hconfig][3] [7]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][3] [7]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][3] [7]),
        .O(\syncrregs.r[hrdatas][7]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][7]_i_25 
       (.I0(\slvo[7][hconfig][3] [7]),
        .I1(\slvo[6][hconfig][3] [7]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][3] [7]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][3] [7]),
        .O(\syncrregs.r[hrdatas][7]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][7]_i_26 
       (.I0(\slvo[3][hconfig][0] [7]),
        .I1(\slvo[2][hconfig][0] [7]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][0] [7]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][0] [7]),
        .O(\syncrregs.r[hrdatas][7]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][7]_i_27 
       (.I0(\slvo[7][hconfig][0] [7]),
        .I1(\slvo[6][hconfig][0] [7]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][0] [7]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][0] [7]),
        .O(\syncrregs.r[hrdatas][7]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][7]_i_28 
       (.I0(\slvo[3][hconfig][1] [7]),
        .I1(\slvo[2][hconfig][1] [7]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][1] [7]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][1] [7]),
        .O(\syncrregs.r[hrdatas][7]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][7]_i_29 
       (.I0(\slvo[7][hconfig][1] [7]),
        .I1(\slvo[6][hconfig][1] [7]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][1] [7]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][1] [7]),
        .O(\syncrregs.r[hrdatas][7]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][8]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][8]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][8]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][8]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][8]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][8]_i_14 
       (.I0(\slvo[3][hconfig][6] [8]),
        .I1(\slvo[2][hconfig][6] [8]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][6] [8]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][6] [8]),
        .O(\syncrregs.r[hrdatas][8]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][8]_i_15 
       (.I0(\slvo[7][hconfig][6] [8]),
        .I1(\slvo[6][hconfig][6] [8]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][6] [8]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][6] [8]),
        .O(\syncrregs.r[hrdatas][8]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][8]_i_16 
       (.I0(\slvo[3][hconfig][7] [8]),
        .I1(\slvo[2][hconfig][7] [8]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][7] [8]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][7] [8]),
        .O(\syncrregs.r[hrdatas][8]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][8]_i_17 
       (.I0(\slvo[7][hconfig][7] [8]),
        .I1(\slvo[6][hconfig][7] [8]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][7] [8]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][7] [8]),
        .O(\syncrregs.r[hrdatas][8]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][8]_i_18 
       (.I0(\slvo[3][hconfig][4] [8]),
        .I1(\slvo[2][hconfig][4] [8]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][4] [8]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][4] [8]),
        .O(\syncrregs.r[hrdatas][8]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][8]_i_19 
       (.I0(\slvo[7][hconfig][4] [8]),
        .I1(\slvo[6][hconfig][4] [8]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][4] [8]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][4] [8]),
        .O(\syncrregs.r[hrdatas][8]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][8]_i_20 
       (.I0(\slvo[3][hconfig][5] [8]),
        .I1(\slvo[2][hconfig][5] [8]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][5] [8]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][5] [8]),
        .O(\syncrregs.r[hrdatas][8]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][8]_i_21 
       (.I0(\slvo[7][hconfig][5] [8]),
        .I1(\slvo[6][hconfig][5] [8]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][5] [8]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][5] [8]),
        .O(\syncrregs.r[hrdatas][8]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][8]_i_22 
       (.I0(\slvo[3][hconfig][2] [8]),
        .I1(\slvo[2][hconfig][2] [8]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][2] [8]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][2] [8]),
        .O(\syncrregs.r[hrdatas][8]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][8]_i_23 
       (.I0(\slvo[7][hconfig][2] [8]),
        .I1(\slvo[6][hconfig][2] [8]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][2] [8]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][2] [8]),
        .O(\syncrregs.r[hrdatas][8]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][8]_i_24 
       (.I0(\slvo[3][hconfig][3] [8]),
        .I1(\slvo[2][hconfig][3] [8]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][3] [8]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][3] [8]),
        .O(\syncrregs.r[hrdatas][8]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][8]_i_25 
       (.I0(\slvo[7][hconfig][3] [8]),
        .I1(\slvo[6][hconfig][3] [8]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][3] [8]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][3] [8]),
        .O(\syncrregs.r[hrdatas][8]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][8]_i_26 
       (.I0(\slvo[3][hconfig][0] [8]),
        .I1(\slvo[2][hconfig][0] [8]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][0] [8]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][0] [8]),
        .O(\syncrregs.r[hrdatas][8]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][8]_i_27 
       (.I0(\slvo[7][hconfig][0] [8]),
        .I1(\slvo[6][hconfig][0] [8]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][0] [8]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][0] [8]),
        .O(\syncrregs.r[hrdatas][8]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][8]_i_28 
       (.I0(\slvo[3][hconfig][1] [8]),
        .I1(\slvo[2][hconfig][1] [8]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][1] [8]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][1] [8]),
        .O(\syncrregs.r[hrdatas][8]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][8]_i_29 
       (.I0(\slvo[7][hconfig][1] [8]),
        .I1(\slvo[6][hconfig][1] [8]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][1] [8]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][1] [8]),
        .O(\syncrregs.r[hrdatas][8]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][9]_i_1 
       (.I0(\syncrregs.r_reg[hrdatas][9]_i_2_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][9]_i_3_n_0 ),
        .I2(\syncrregs.r_reg[haddr_n_0_][4] ),
        .I3(\syncrregs.r_reg[hrdatas][9]_i_4_n_0 ),
        .I4(\syncrregs.r_reg[haddr_n_0_][3] ),
        .I5(\syncrregs.r_reg[hrdatas][9]_i_5_n_0 ),
        .O(\slvo[15][hready]__0 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][9]_i_14 
       (.I0(\slvo[3][hconfig][6] [9]),
        .I1(\slvo[2][hconfig][6] [9]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][6] [9]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][6] [9]),
        .O(\syncrregs.r[hrdatas][9]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][9]_i_15 
       (.I0(\slvo[7][hconfig][6] [9]),
        .I1(\slvo[6][hconfig][6] [9]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][6] [9]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][6] [9]),
        .O(\syncrregs.r[hrdatas][9]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][9]_i_16 
       (.I0(\slvo[3][hconfig][7] [9]),
        .I1(\slvo[2][hconfig][7] [9]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][7] [9]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][7] [9]),
        .O(\syncrregs.r[hrdatas][9]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][9]_i_17 
       (.I0(\slvo[7][hconfig][7] [9]),
        .I1(\slvo[6][hconfig][7] [9]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][7] [9]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][7] [9]),
        .O(\syncrregs.r[hrdatas][9]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][9]_i_18 
       (.I0(\slvo[3][hconfig][4] [9]),
        .I1(\slvo[2][hconfig][4] [9]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][4] [9]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][4] [9]),
        .O(\syncrregs.r[hrdatas][9]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][9]_i_19 
       (.I0(\slvo[7][hconfig][4] [9]),
        .I1(\slvo[6][hconfig][4] [9]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][4] [9]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][4] [9]),
        .O(\syncrregs.r[hrdatas][9]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][9]_i_20 
       (.I0(\slvo[3][hconfig][5] [9]),
        .I1(\slvo[2][hconfig][5] [9]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][5] [9]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][5] [9]),
        .O(\syncrregs.r[hrdatas][9]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][9]_i_21 
       (.I0(\slvo[7][hconfig][5] [9]),
        .I1(\slvo[6][hconfig][5] [9]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][5] [9]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][5] [9]),
        .O(\syncrregs.r[hrdatas][9]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][9]_i_22 
       (.I0(\slvo[3][hconfig][2] [9]),
        .I1(\slvo[2][hconfig][2] [9]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][2] [9]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][2] [9]),
        .O(\syncrregs.r[hrdatas][9]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][9]_i_23 
       (.I0(\slvo[7][hconfig][2] [9]),
        .I1(\slvo[6][hconfig][2] [9]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][2] [9]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][2] [9]),
        .O(\syncrregs.r[hrdatas][9]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][9]_i_24 
       (.I0(\slvo[3][hconfig][3] [9]),
        .I1(\slvo[2][hconfig][3] [9]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][3] [9]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][3] [9]),
        .O(\syncrregs.r[hrdatas][9]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][9]_i_25 
       (.I0(\slvo[7][hconfig][3] [9]),
        .I1(\slvo[6][hconfig][3] [9]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][3] [9]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][3] [9]),
        .O(\syncrregs.r[hrdatas][9]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][9]_i_26 
       (.I0(\slvo[3][hconfig][0] [9]),
        .I1(\slvo[2][hconfig][0] [9]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][0] [9]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][0] [9]),
        .O(\syncrregs.r[hrdatas][9]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][9]_i_27 
       (.I0(\slvo[7][hconfig][0] [9]),
        .I1(\slvo[6][hconfig][0] [9]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][0] [9]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][0] [9]),
        .O(\syncrregs.r[hrdatas][9]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][9]_i_28 
       (.I0(\slvo[3][hconfig][1] [9]),
        .I1(\slvo[2][hconfig][1] [9]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[1][hconfig][1] [9]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[0][hconfig][1] [9]),
        .O(\syncrregs.r[hrdatas][9]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \syncrregs.r[hrdatas][9]_i_29 
       (.I0(\slvo[7][hconfig][1] [9]),
        .I1(\slvo[6][hconfig][1] [9]),
        .I2(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .I3(\slvo[5][hconfig][1] [9]),
        .I4(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .I5(\slvo[4][hconfig][1] [9]),
        .O(\syncrregs.r[hrdatas][9]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0E00)) 
    \syncrregs.r[hready]_i_1 
       (.I0(\syncrregs.r_reg[defslv]__0 ),
        .I1(\syncrregs.r_reg[cfgsel_n_0_] ),
        .I2(\syncrregs.r_reg[hready_n_0_] ),
        .I3(\syncrregs.r_reg[htrans_n_0_][1] ),
        .O(rin));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \syncrregs.r[hslave][0]_i_1 
       (.I0(\slvi[hsel][7]_INST_0_i_1_n_0 ),
        .I1(\slvi[hsel][1]_INST_0_i_1_n_0 ),
        .I2(p_0_in5_in),
        .I3(p_2_in),
        .O(p_6_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \syncrregs.r[hslave][1]_i_1 
       (.I0(p_0_in5_in),
        .I1(\slvi[hsel][7]_INST_0_i_1_n_0 ),
        .I2(p_1_in10_in),
        .I3(p_2_in7_in),
        .O(p_11_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \syncrregs.r[hslave][2]_i_1 
       (.I0(p_2_in),
        .I1(\slvi[hsel][7]_INST_0_i_1_n_0 ),
        .I2(p_2_in7_in),
        .I3(p_1_in13_in),
        .O(p_14_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \syncrregs.r[htrans][1]_i_1 
       (.I0(rst),
        .O(\syncrregs.r[htrans][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[cfga11] 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\slvi[haddr] [11]),
        .Q(\syncrregs.r_reg ),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[cfgsel] 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(hsel1192_out),
        .Q(\syncrregs.r_reg[cfgsel_n_0_] ),
        .R(\syncrregs.r[htrans][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[defslv] 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(p_185_out),
        .Q(\syncrregs.r_reg[defslv]__0 ),
        .R(\syncrregs.r[htrans][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[haddr][10] 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\slvi[haddr] [10]),
        .Q(sel0[6]),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[haddr][2] 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\slvi[haddr] [2]),
        .Q(\syncrregs.r_reg[haddr_n_0_][2] ),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[haddr][3] 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\slvi[haddr] [3]),
        .Q(\syncrregs.r_reg[haddr_n_0_][3] ),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[haddr][4] 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\slvi[haddr] [4]),
        .Q(\syncrregs.r_reg[haddr_n_0_][4] ),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "syncrregs.r_reg[haddr][5]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[haddr][5] 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\slvi[haddr] [5]),
        .Q(sel0[1]),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "syncrregs.r_reg[haddr][5]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[haddr][5]_rep 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\slvi[haddr] [5]),
        .Q(\syncrregs.r_reg[haddr][5]_rep_n_0 ),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "syncrregs.r_reg[haddr][5]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[haddr][5]_rep__0 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\slvi[haddr] [5]),
        .Q(\syncrregs.r_reg[haddr][5]_rep__0_n_0 ),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "syncrregs.r_reg[haddr][5]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[haddr][5]_rep__1 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\slvi[haddr] [5]),
        .Q(\syncrregs.r_reg[haddr][5]_rep__1_n_0 ),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "syncrregs.r_reg[haddr][5]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[haddr][5]_rep__2 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\slvi[haddr] [5]),
        .Q(\syncrregs.r_reg[haddr][5]_rep__2_n_0 ),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "syncrregs.r_reg[haddr][5]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[haddr][5]_rep__3 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\slvi[haddr] [5]),
        .Q(\syncrregs.r_reg[haddr][5]_rep__3_n_0 ),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "syncrregs.r_reg[haddr][6]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[haddr][6] 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\slvi[haddr] [6]),
        .Q(sel0[2]),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "syncrregs.r_reg[haddr][6]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[haddr][6]_rep 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\slvi[haddr] [6]),
        .Q(\syncrregs.r_reg[haddr][6]_rep_n_0 ),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "syncrregs.r_reg[haddr][6]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[haddr][6]_rep__0 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\slvi[haddr] [6]),
        .Q(\syncrregs.r_reg[haddr][6]_rep__0_n_0 ),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "syncrregs.r_reg[haddr][6]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[haddr][6]_rep__1 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\slvi[haddr] [6]),
        .Q(\syncrregs.r_reg[haddr][6]_rep__1_n_0 ),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "syncrregs.r_reg[haddr][6]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[haddr][6]_rep__2 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\slvi[haddr] [6]),
        .Q(\syncrregs.r_reg[haddr][6]_rep__2_n_0 ),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "syncrregs.r_reg[haddr][6]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[haddr][6]_rep__3 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\slvi[haddr] [6]),
        .Q(\syncrregs.r_reg[haddr][6]_rep__3_n_0 ),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "syncrregs.r_reg[haddr][7]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[haddr][7] 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\slvi[haddr] [7]),
        .Q(sel0[3]),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "syncrregs.r_reg[haddr][7]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[haddr][7]_rep 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\slvi[haddr] [7]),
        .Q(\syncrregs.r_reg[haddr][7]_rep_n_0 ),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "syncrregs.r_reg[haddr][7]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[haddr][7]_rep__0 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\slvi[haddr] [7]),
        .Q(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[haddr][8] 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\slvi[haddr] [8]),
        .Q(sel0[4]),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[haddr][9] 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\slvi[haddr] [9]),
        .Q(sel0[5]),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hmaster][0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r ),
        .Q(\^slvi[hmaster] [0]),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hmaster][1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r[hmaster][1]_i_1_n_0 ),
        .Q(\^slvi[hmaster] [1]),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hmaster][2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r[hmaster][2]_i_1_n_0 ),
        .Q(\^slvi[hmaster] [2]),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hmasterd][0] 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\^slvi[hmaster] [0]),
        .Q(\syncrregs.r_reg[hmasterd]__0 [0]),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hmasterd][1] 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\^slvi[hmaster] [1]),
        .Q(\syncrregs.r_reg[hmasterd]__0 [1]),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hmasterd][2] 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\^slvi[hmaster] [2]),
        .Q(\syncrregs.r_reg[hmasterd]__0 [2]),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hmasterlock] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r[hmasterlock]_i_1_n_0 ),
        .Q(\slvi[hmastlock] ),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hmasterlock]_i_2 
       (.I0(\syncrregs.r[hmasterlock]_i_4_n_0 ),
        .I1(\syncrregs.r[hmasterlock]_i_5_n_0 ),
        .O(\syncrregs.r_reg[hmasterlock]_i_2_n_0 ),
        .S(\syncrregs.r[hmaster][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hmasterlockd] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r[hmasterlockd]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hmasterlockd]__0 ),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][0]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [0]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][0]_i_1 
       (.I0(\syncrregs.r[hrdatam][0]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][0]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][0]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][10]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [10]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][10]_i_1 
       (.I0(\syncrregs.r[hrdatam][10]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][10]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][10]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][11]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [11]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][11]_i_1 
       (.I0(\syncrregs.r[hrdatam][11]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][11]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][11]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][12]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [12]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][12]_i_1 
       (.I0(\syncrregs.r[hrdatam][12]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][12]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][12]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][13]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [13]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][13]_i_1 
       (.I0(\syncrregs.r[hrdatam][13]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][13]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][13]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][14]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [14]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][14]_i_1 
       (.I0(\syncrregs.r[hrdatam][14]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][14]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][14]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][15]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [15]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][15]_i_1 
       (.I0(\syncrregs.r[hrdatam][15]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][15]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][15]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][16]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [16]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][16]_i_1 
       (.I0(\syncrregs.r[hrdatam][16]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][16]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][16]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][17]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [17]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][17]_i_1 
       (.I0(\syncrregs.r[hrdatam][17]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][17]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][17]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][18]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [18]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][18]_i_1 
       (.I0(\syncrregs.r[hrdatam][18]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][18]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][18]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][19]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [19]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][19]_i_1 
       (.I0(\syncrregs.r[hrdatam][19]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][19]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][19]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][1]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [1]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][1]_i_1 
       (.I0(\syncrregs.r[hrdatam][1]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][1]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][1]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][20]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [20]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][20]_i_1 
       (.I0(\syncrregs.r[hrdatam][20]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][20]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][20]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][21]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [21]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][21]_i_1 
       (.I0(\syncrregs.r[hrdatam][21]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][21]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][21]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][22]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [22]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][22]_i_1 
       (.I0(\syncrregs.r[hrdatam][22]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][22]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][22]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][23]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [23]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][23]_i_1 
       (.I0(\syncrregs.r[hrdatam][23]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][23]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][23]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][24]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [24]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][24]_i_1 
       (.I0(\syncrregs.r[hrdatam][24]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][24]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][24]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][25]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [25]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][25]_i_1 
       (.I0(\syncrregs.r[hrdatam][25]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][25]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][25]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][26]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [26]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][26]_i_1 
       (.I0(\syncrregs.r[hrdatam][26]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][26]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][26]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][27]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [27]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][27]_i_1 
       (.I0(\syncrregs.r[hrdatam][27]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][27]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][27]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][28]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [28]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][28]_i_1 
       (.I0(\syncrregs.r[hrdatam][28]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][28]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][28]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][29]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [29]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][29]_i_1 
       (.I0(\syncrregs.r[hrdatam][29]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][29]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][29]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][2]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [2]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][2]_i_1 
       (.I0(\syncrregs.r[hrdatam][2]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][2]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][2]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][30]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [30]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][30]_i_1 
       (.I0(\syncrregs.r[hrdatam][30]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][30]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][30]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][31]_i_2_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [31]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][31]_i_2 
       (.I0(\syncrregs.r[hrdatam][31]_i_3_n_0 ),
        .I1(\syncrregs.r[hrdatam][31]_i_4_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][31]_i_2_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][3]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [3]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][3]_i_1 
       (.I0(\syncrregs.r[hrdatam][3]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][3]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][3]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][4]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [4]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][4]_i_1 
       (.I0(\syncrregs.r[hrdatam][4]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][4]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][4]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][5]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [5]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][5]_i_1 
       (.I0(\syncrregs.r[hrdatam][5]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][5]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][5]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][6]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [6]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][6]_i_1 
       (.I0(\syncrregs.r[hrdatam][6]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][6]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][6]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][7]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [7]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][7]_i_1 
       (.I0(\syncrregs.r[hrdatam][7]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][7]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][7]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][8]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [8]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][8]_i_1 
       (.I0(\syncrregs.r[hrdatam][8]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][8]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][8]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatam][9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r_reg[hrdatam][9]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatam]__0 [9]),
        .R(\syncrregs.r[hrdatam][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatam][9]_i_1 
       (.I0(\syncrregs.r[hrdatam][9]_i_2_n_0 ),
        .I1(\syncrregs.r[hrdatam][9]_i_3_n_0 ),
        .O(\syncrregs.r_reg[hrdatam][9]_i_1_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [0]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [0]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][0]_i_10 
       (.I0(\syncrregs.r[hrdatas][0]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][0]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][0]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][0]_i_11 
       (.I0(\syncrregs.r[hrdatas][0]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][0]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][0]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][0]_i_12 
       (.I0(\syncrregs.r[hrdatas][0]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][0]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][0]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][0]_i_13 
       (.I0(\syncrregs.r[hrdatas][0]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][0]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][0]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][0]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][0]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][0]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][0]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][0]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][0]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][0]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][0]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][0]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][0]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][0]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][0]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][0]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][0]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][0]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][0]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][0]_i_6 
       (.I0(\syncrregs.r[hrdatas][0]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][0]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][0]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][0]_i_7 
       (.I0(\syncrregs.r[hrdatas][0]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][0]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][0]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][0]_i_8 
       (.I0(\syncrregs.r[hrdatas][0]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][0]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][0]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][0]_i_9 
       (.I0(\syncrregs.r[hrdatas][0]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][0]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][0]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [10]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [10]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][10]_i_10 
       (.I0(\syncrregs.r[hrdatas][10]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][10]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][10]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][10]_i_11 
       (.I0(\syncrregs.r[hrdatas][10]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][10]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][10]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][10]_i_12 
       (.I0(\syncrregs.r[hrdatas][10]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][10]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][10]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][10]_i_13 
       (.I0(\syncrregs.r[hrdatas][10]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][10]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][10]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][10]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][10]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][10]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][10]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][10]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][10]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][10]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][10]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][10]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][10]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][10]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][10]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][10]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][10]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][10]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][10]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][10]_i_6 
       (.I0(\syncrregs.r[hrdatas][10]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][10]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][10]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][10]_i_7 
       (.I0(\syncrregs.r[hrdatas][10]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][10]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][10]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][10]_i_8 
       (.I0(\syncrregs.r[hrdatas][10]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][10]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][10]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][10]_i_9 
       (.I0(\syncrregs.r[hrdatas][10]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][10]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][10]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [11]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [11]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][11]_i_10 
       (.I0(\syncrregs.r[hrdatas][11]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][11]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][11]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][11]_i_11 
       (.I0(\syncrregs.r[hrdatas][11]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][11]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][11]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][11]_i_12 
       (.I0(\syncrregs.r[hrdatas][11]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][11]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][11]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][11]_i_13 
       (.I0(\syncrregs.r[hrdatas][11]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][11]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][11]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][11]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][11]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][11]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][11]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][11]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][11]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][11]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][11]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][11]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][11]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][11]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][11]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][11]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][11]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][11]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][11]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][11]_i_6 
       (.I0(\syncrregs.r[hrdatas][11]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][11]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][11]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][11]_i_7 
       (.I0(\syncrregs.r[hrdatas][11]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][11]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][11]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][11]_i_8 
       (.I0(\syncrregs.r[hrdatas][11]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][11]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][11]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][11]_i_9 
       (.I0(\syncrregs.r[hrdatas][11]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][11]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][11]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r[hrdatas][12]_i_2_n_0 ),
        .Q(\syncrregs.r_reg[hrdatas]__0 [12]),
        .S(\v[hrdatas] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][12]_i_10 
       (.I0(\syncrregs.r[hrdatas][12]_i_21_n_0 ),
        .I1(\syncrregs.r[hrdatas][12]_i_22_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][12]_i_10_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][12]_i_11 
       (.I0(\syncrregs.r[hrdatas][12]_i_23_n_0 ),
        .I1(\syncrregs.r[hrdatas][12]_i_24_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][12]_i_11_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][12]_i_12 
       (.I0(\syncrregs.r[hrdatas][12]_i_25_n_0 ),
        .I1(\syncrregs.r[hrdatas][12]_i_26_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][12]_i_12_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][12]_i_13 
       (.I0(\syncrregs.r[hrdatas][12]_i_27_n_0 ),
        .I1(\syncrregs.r[hrdatas][12]_i_28_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][12]_i_13_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][12]_i_14 
       (.I0(\syncrregs.r[hrdatas][12]_i_29_n_0 ),
        .I1(\syncrregs.r[hrdatas][12]_i_30_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][12]_i_14_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][12]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][12]_i_11_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][12]_i_12_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][12]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][12]_i_6 
       (.I0(\syncrregs.r_reg[hrdatas][12]_i_13_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][12]_i_14_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][12]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][12]_i_7 
       (.I0(\syncrregs.r[hrdatas][12]_i_15_n_0 ),
        .I1(\syncrregs.r[hrdatas][12]_i_16_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][12]_i_7_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][12]_i_8 
       (.I0(\syncrregs.r[hrdatas][12]_i_17_n_0 ),
        .I1(\syncrregs.r[hrdatas][12]_i_18_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][12]_i_8_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][12]_i_9 
       (.I0(\syncrregs.r[hrdatas][12]_i_19_n_0 ),
        .I1(\syncrregs.r[hrdatas][12]_i_20_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][12]_i_9_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [13]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [13]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][13]_i_10 
       (.I0(\syncrregs.r[hrdatas][13]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][13]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][13]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][13]_i_11 
       (.I0(\syncrregs.r[hrdatas][13]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][13]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][13]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][13]_i_12 
       (.I0(\syncrregs.r[hrdatas][13]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][13]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][13]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][13]_i_13 
       (.I0(\syncrregs.r[hrdatas][13]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][13]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][13]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][13]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][13]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][13]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][13]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][13]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][13]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][13]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][13]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][13]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][13]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][13]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][13]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][13]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][13]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][13]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][13]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][13]_i_6 
       (.I0(\syncrregs.r[hrdatas][13]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][13]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][13]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][13]_i_7 
       (.I0(\syncrregs.r[hrdatas][13]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][13]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][13]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][13]_i_8 
       (.I0(\syncrregs.r[hrdatas][13]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][13]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][13]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][13]_i_9 
       (.I0(\syncrregs.r[hrdatas][13]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][13]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][13]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [14]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [14]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][14]_i_10 
       (.I0(\syncrregs.r[hrdatas][14]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][14]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][14]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][14]_i_11 
       (.I0(\syncrregs.r[hrdatas][14]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][14]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][14]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][14]_i_12 
       (.I0(\syncrregs.r[hrdatas][14]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][14]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][14]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][14]_i_13 
       (.I0(\syncrregs.r[hrdatas][14]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][14]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][14]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][14]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][14]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][14]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][14]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][14]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][14]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][14]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][14]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][14]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][14]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][14]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][14]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][14]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][14]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][14]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][14]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][14]_i_6 
       (.I0(\syncrregs.r[hrdatas][14]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][14]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][14]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][14]_i_7 
       (.I0(\syncrregs.r[hrdatas][14]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][14]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][14]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][14]_i_8 
       (.I0(\syncrregs.r[hrdatas][14]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][14]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][14]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][14]_i_9 
       (.I0(\syncrregs.r[hrdatas][14]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][14]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][14]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [15]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [15]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][15]_i_10 
       (.I0(\syncrregs.r[hrdatas][15]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][15]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][15]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][15]_i_11 
       (.I0(\syncrregs.r[hrdatas][15]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][15]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][15]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][15]_i_12 
       (.I0(\syncrregs.r[hrdatas][15]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][15]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][15]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][15]_i_13 
       (.I0(\syncrregs.r[hrdatas][15]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][15]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][15]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][15]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][15]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][15]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][15]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][15]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][15]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][15]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][15]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][15]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][15]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][15]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][15]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][15]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][15]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][15]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][15]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][15]_i_6 
       (.I0(\syncrregs.r[hrdatas][15]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][15]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][15]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][15]_i_7 
       (.I0(\syncrregs.r[hrdatas][15]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][15]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][15]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][15]_i_8 
       (.I0(\syncrregs.r[hrdatas][15]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][15]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][15]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][15]_i_9 
       (.I0(\syncrregs.r[hrdatas][15]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][15]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][15]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [16]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [16]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][16]_i_10 
       (.I0(\syncrregs.r[hrdatas][16]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][16]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][16]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][16]_i_11 
       (.I0(\syncrregs.r[hrdatas][16]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][16]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][16]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][16]_i_12 
       (.I0(\syncrregs.r[hrdatas][16]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][16]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][16]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][16]_i_13 
       (.I0(\syncrregs.r[hrdatas][16]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][16]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][16]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][16]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][16]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][16]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][16]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][16]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][16]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][16]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][16]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][16]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][16]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][16]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][16]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][16]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][16]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][16]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][16]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][16]_i_6 
       (.I0(\syncrregs.r[hrdatas][16]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][16]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][16]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][16]_i_7 
       (.I0(\syncrregs.r[hrdatas][16]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][16]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][16]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][16]_i_8 
       (.I0(\syncrregs.r[hrdatas][16]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][16]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][16]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][16]_i_9 
       (.I0(\syncrregs.r[hrdatas][16]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][16]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][16]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [17]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [17]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][17]_i_10 
       (.I0(\syncrregs.r[hrdatas][17]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][17]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][17]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][17]_i_11 
       (.I0(\syncrregs.r[hrdatas][17]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][17]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][17]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][17]_i_12 
       (.I0(\syncrregs.r[hrdatas][17]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][17]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][17]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][17]_i_13 
       (.I0(\syncrregs.r[hrdatas][17]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][17]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][17]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][17]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][17]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][17]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][17]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][17]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][17]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][17]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][17]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][17]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][17]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][17]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][17]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][17]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][17]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][17]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][17]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][17]_i_6 
       (.I0(\syncrregs.r[hrdatas][17]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][17]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][17]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][17]_i_7 
       (.I0(\syncrregs.r[hrdatas][17]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][17]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][17]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][17]_i_8 
       (.I0(\syncrregs.r[hrdatas][17]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][17]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][17]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][17]_i_9 
       (.I0(\syncrregs.r[hrdatas][17]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][17]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][17]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [18]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [18]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][18]_i_10 
       (.I0(\syncrregs.r[hrdatas][18]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][18]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][18]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][18]_i_11 
       (.I0(\syncrregs.r[hrdatas][18]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][18]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][18]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][18]_i_12 
       (.I0(\syncrregs.r[hrdatas][18]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][18]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][18]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][18]_i_13 
       (.I0(\syncrregs.r[hrdatas][18]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][18]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][18]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][18]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][18]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][18]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][18]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][18]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][18]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][18]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][18]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][18]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][18]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][18]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][18]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][18]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][18]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][18]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][18]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][18]_i_6 
       (.I0(\syncrregs.r[hrdatas][18]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][18]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][18]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][18]_i_7 
       (.I0(\syncrregs.r[hrdatas][18]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][18]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][18]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][18]_i_8 
       (.I0(\syncrregs.r[hrdatas][18]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][18]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][18]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][18]_i_9 
       (.I0(\syncrregs.r[hrdatas][18]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][18]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][18]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [19]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [19]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][19]_i_10 
       (.I0(\syncrregs.r[hrdatas][19]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][19]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][19]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][19]_i_11 
       (.I0(\syncrregs.r[hrdatas][19]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][19]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][19]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][19]_i_12 
       (.I0(\syncrregs.r[hrdatas][19]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][19]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][19]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][19]_i_13 
       (.I0(\syncrregs.r[hrdatas][19]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][19]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][19]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][19]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][19]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][19]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][19]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][19]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][19]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][19]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][19]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][19]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][19]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][19]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][19]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][19]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][19]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][19]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][19]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][19]_i_6 
       (.I0(\syncrregs.r[hrdatas][19]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][19]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][19]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][19]_i_7 
       (.I0(\syncrregs.r[hrdatas][19]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][19]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][19]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][19]_i_8 
       (.I0(\syncrregs.r[hrdatas][19]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][19]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][19]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][19]_i_9 
       (.I0(\syncrregs.r[hrdatas][19]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][19]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][19]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r[hrdatas][1]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatas]__0 [1]),
        .S(\v[hrdatas] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][1]_i_10 
       (.I0(\syncrregs.r[hrdatas][1]_i_23_n_0 ),
        .I1(\syncrregs.r[hrdatas][1]_i_24_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][1]_i_10_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][1]_i_11 
       (.I0(\syncrregs.r[hrdatas][1]_i_25_n_0 ),
        .I1(\syncrregs.r[hrdatas][1]_i_26_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][1]_i_11_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][1]_i_12 
       (.I0(\syncrregs.r[hrdatas][1]_i_27_n_0 ),
        .I1(\syncrregs.r[hrdatas][1]_i_28_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][1]_i_12_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][1]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][1]_i_9_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][1]_i_10_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][1]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][1]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][1]_i_11_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][1]_i_12_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][1]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][1]_i_5 
       (.I0(\syncrregs.r[hrdatas][1]_i_13_n_0 ),
        .I1(\syncrregs.r[hrdatas][1]_i_14_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][1]_i_5_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][1]_i_6 
       (.I0(\syncrregs.r[hrdatas][1]_i_15_n_0 ),
        .I1(\syncrregs.r[hrdatas][1]_i_16_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][1]_i_6_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][1]_i_7 
       (.I0(\syncrregs.r[hrdatas][1]_i_17_n_0 ),
        .I1(\syncrregs.r[hrdatas][1]_i_18_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][1]_i_7_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][1]_i_8 
       (.I0(\syncrregs.r[hrdatas][1]_i_19_n_0 ),
        .I1(\syncrregs.r[hrdatas][1]_i_20_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][1]_i_8_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][1]_i_9 
       (.I0(\syncrregs.r[hrdatas][1]_i_21_n_0 ),
        .I1(\syncrregs.r[hrdatas][1]_i_22_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][1]_i_9_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [20]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [20]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][20]_i_10 
       (.I0(\syncrregs.r[hrdatas][20]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][20]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][20]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][20]_i_11 
       (.I0(\syncrregs.r[hrdatas][20]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][20]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][20]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][20]_i_12 
       (.I0(\syncrregs.r[hrdatas][20]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][20]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][20]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][20]_i_13 
       (.I0(\syncrregs.r[hrdatas][20]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][20]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][20]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][20]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][20]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][20]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][20]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][20]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][20]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][20]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][20]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][20]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][20]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][20]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][20]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][20]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][20]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][20]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][20]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][20]_i_6 
       (.I0(\syncrregs.r[hrdatas][20]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][20]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][20]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][20]_i_7 
       (.I0(\syncrregs.r[hrdatas][20]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][20]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][20]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][20]_i_8 
       (.I0(\syncrregs.r[hrdatas][20]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][20]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][20]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][20]_i_9 
       (.I0(\syncrregs.r[hrdatas][20]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][20]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][20]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [21]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [21]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][21]_i_10 
       (.I0(\syncrregs.r[hrdatas][21]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][21]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][21]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][21]_i_11 
       (.I0(\syncrregs.r[hrdatas][21]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][21]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][21]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][21]_i_12 
       (.I0(\syncrregs.r[hrdatas][21]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][21]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][21]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][21]_i_13 
       (.I0(\syncrregs.r[hrdatas][21]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][21]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][21]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][21]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][21]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][21]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][21]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][21]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][21]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][21]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][21]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][21]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][21]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][21]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][21]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][21]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][21]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][21]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][21]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][21]_i_6 
       (.I0(\syncrregs.r[hrdatas][21]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][21]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][21]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][21]_i_7 
       (.I0(\syncrregs.r[hrdatas][21]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][21]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][21]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][21]_i_8 
       (.I0(\syncrregs.r[hrdatas][21]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][21]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][21]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][21]_i_9 
       (.I0(\syncrregs.r[hrdatas][21]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][21]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][21]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [22]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [22]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][22]_i_10 
       (.I0(\syncrregs.r[hrdatas][22]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][22]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][22]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][22]_i_11 
       (.I0(\syncrregs.r[hrdatas][22]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][22]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][22]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][22]_i_12 
       (.I0(\syncrregs.r[hrdatas][22]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][22]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][22]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][22]_i_13 
       (.I0(\syncrregs.r[hrdatas][22]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][22]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][22]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][22]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][22]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][22]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][22]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][22]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][22]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][22]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][22]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][22]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][22]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][22]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][22]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][22]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][22]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][22]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][22]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][22]_i_6 
       (.I0(\syncrregs.r[hrdatas][22]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][22]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][22]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][22]_i_7 
       (.I0(\syncrregs.r[hrdatas][22]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][22]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][22]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][22]_i_8 
       (.I0(\syncrregs.r[hrdatas][22]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][22]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][22]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][22]_i_9 
       (.I0(\syncrregs.r[hrdatas][22]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][22]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][22]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [23]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [23]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][23]_i_10 
       (.I0(\syncrregs.r[hrdatas][23]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][23]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][23]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][23]_i_11 
       (.I0(\syncrregs.r[hrdatas][23]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][23]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][23]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][23]_i_12 
       (.I0(\syncrregs.r[hrdatas][23]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][23]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][23]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][23]_i_13 
       (.I0(\syncrregs.r[hrdatas][23]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][23]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][23]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][23]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][23]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][23]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][23]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][23]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][23]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][23]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][23]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][23]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][23]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][23]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][23]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][23]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][23]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][23]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][23]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][23]_i_6 
       (.I0(\syncrregs.r[hrdatas][23]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][23]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][23]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][23]_i_7 
       (.I0(\syncrregs.r[hrdatas][23]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][23]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][23]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][23]_i_8 
       (.I0(\syncrregs.r[hrdatas][23]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][23]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][23]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][23]_i_9 
       (.I0(\syncrregs.r[hrdatas][23]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][23]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][23]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [24]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [24]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][24]_i_10 
       (.I0(\syncrregs.r[hrdatas][24]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][24]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][24]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][24]_i_11 
       (.I0(\syncrregs.r[hrdatas][24]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][24]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][24]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][24]_i_12 
       (.I0(\syncrregs.r[hrdatas][24]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][24]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][24]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][24]_i_13 
       (.I0(\syncrregs.r[hrdatas][24]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][24]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][24]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][24]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][24]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][24]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][24]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][24]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][24]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][24]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][24]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][24]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][24]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][24]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][24]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][24]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][24]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][24]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][24]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][24]_i_6 
       (.I0(\syncrregs.r[hrdatas][24]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][24]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][24]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][24]_i_7 
       (.I0(\syncrregs.r[hrdatas][24]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][24]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][24]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][24]_i_8 
       (.I0(\syncrregs.r[hrdatas][24]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][24]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][24]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][24]_i_9 
       (.I0(\syncrregs.r[hrdatas][24]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][24]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][24]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [25]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [25]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][25]_i_10 
       (.I0(\syncrregs.r[hrdatas][25]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][25]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][25]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][25]_i_11 
       (.I0(\syncrregs.r[hrdatas][25]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][25]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][25]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][25]_i_12 
       (.I0(\syncrregs.r[hrdatas][25]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][25]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][25]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][25]_i_13 
       (.I0(\syncrregs.r[hrdatas][25]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][25]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][25]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][25]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][25]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][25]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][25]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][25]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][25]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][25]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][25]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][25]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][25]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][25]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][25]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][25]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][25]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][25]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][25]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][25]_i_6 
       (.I0(\syncrregs.r[hrdatas][25]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][25]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][25]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][25]_i_7 
       (.I0(\syncrregs.r[hrdatas][25]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][25]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][25]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][25]_i_8 
       (.I0(\syncrregs.r[hrdatas][25]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][25]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][25]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][25]_i_9 
       (.I0(\syncrregs.r[hrdatas][25]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][25]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][25]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [26]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [26]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][26]_i_10 
       (.I0(\syncrregs.r[hrdatas][26]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][26]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][26]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][26]_i_11 
       (.I0(\syncrregs.r[hrdatas][26]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][26]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][26]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][26]_i_12 
       (.I0(\syncrregs.r[hrdatas][26]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][26]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][26]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][26]_i_13 
       (.I0(\syncrregs.r[hrdatas][26]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][26]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][26]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][26]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][26]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][26]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][26]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][26]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][26]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][26]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][26]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][26]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][26]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][26]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][26]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][26]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][26]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][26]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][26]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][26]_i_6 
       (.I0(\syncrregs.r[hrdatas][26]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][26]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][26]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][26]_i_7 
       (.I0(\syncrregs.r[hrdatas][26]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][26]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][26]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][26]_i_8 
       (.I0(\syncrregs.r[hrdatas][26]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][26]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][26]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][26]_i_9 
       (.I0(\syncrregs.r[hrdatas][26]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][26]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][26]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [27]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [27]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][27]_i_10 
       (.I0(\syncrregs.r[hrdatas][27]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][27]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][27]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][27]_i_11 
       (.I0(\syncrregs.r[hrdatas][27]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][27]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][27]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][27]_i_12 
       (.I0(\syncrregs.r[hrdatas][27]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][27]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][27]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][27]_i_13 
       (.I0(\syncrregs.r[hrdatas][27]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][27]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][27]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][27]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][27]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][27]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][27]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][27]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][27]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][27]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][27]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][27]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][27]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][27]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][27]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][27]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][27]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][27]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][27]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][27]_i_6 
       (.I0(\syncrregs.r[hrdatas][27]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][27]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][27]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][27]_i_7 
       (.I0(\syncrregs.r[hrdatas][27]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][27]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][27]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][27]_i_8 
       (.I0(\syncrregs.r[hrdatas][27]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][27]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][27]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][27]_i_9 
       (.I0(\syncrregs.r[hrdatas][27]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][27]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][27]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [28]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [28]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][28]_i_10 
       (.I0(\syncrregs.r[hrdatas][28]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][28]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][28]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][28]_i_11 
       (.I0(\syncrregs.r[hrdatas][28]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][28]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][28]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][28]_i_12 
       (.I0(\syncrregs.r[hrdatas][28]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][28]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][28]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][28]_i_13 
       (.I0(\syncrregs.r[hrdatas][28]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][28]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][28]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][28]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][28]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][28]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][28]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][28]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][28]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][28]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][28]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][28]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][28]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][28]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][28]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][28]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][28]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][28]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][28]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][28]_i_6 
       (.I0(\syncrregs.r[hrdatas][28]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][28]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][28]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][28]_i_7 
       (.I0(\syncrregs.r[hrdatas][28]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][28]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][28]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][28]_i_8 
       (.I0(\syncrregs.r[hrdatas][28]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][28]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][28]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][28]_i_9 
       (.I0(\syncrregs.r[hrdatas][28]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][28]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][28]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [29]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [29]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][29]_i_10 
       (.I0(\syncrregs.r[hrdatas][29]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][29]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][29]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][29]_i_11 
       (.I0(\syncrregs.r[hrdatas][29]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][29]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][29]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][29]_i_12 
       (.I0(\syncrregs.r[hrdatas][29]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][29]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][29]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][29]_i_13 
       (.I0(\syncrregs.r[hrdatas][29]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][29]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][29]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][29]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][29]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][29]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][29]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][29]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][29]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][29]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][29]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][29]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][29]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][29]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][29]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][29]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][29]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][29]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][29]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][29]_i_6 
       (.I0(\syncrregs.r[hrdatas][29]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][29]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][29]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][29]_i_7 
       (.I0(\syncrregs.r[hrdatas][29]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][29]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][29]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][29]_i_8 
       (.I0(\syncrregs.r[hrdatas][29]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][29]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][29]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][29]_i_9 
       (.I0(\syncrregs.r[hrdatas][29]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][29]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][29]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [2]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [2]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][2]_i_10 
       (.I0(\syncrregs.r[hrdatas][2]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][2]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][2]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][2]_i_11 
       (.I0(\syncrregs.r[hrdatas][2]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][2]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][2]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][2]_i_12 
       (.I0(\syncrregs.r[hrdatas][2]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][2]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][2]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][2]_i_13 
       (.I0(\syncrregs.r[hrdatas][2]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][2]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][2]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][2]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][2]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][2]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][2]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][2]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][2]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][2]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][2]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][2]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][2]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][2]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][2]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][2]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][2]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][2]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][2]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][2]_i_6 
       (.I0(\syncrregs.r[hrdatas][2]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][2]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][2]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][2]_i_7 
       (.I0(\syncrregs.r[hrdatas][2]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][2]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][2]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][2]_i_8 
       (.I0(\syncrregs.r[hrdatas][2]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][2]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][2]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][2]_i_9 
       (.I0(\syncrregs.r[hrdatas][2]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][2]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][2]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [30]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [30]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][30]_i_10 
       (.I0(\syncrregs.r[hrdatas][30]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][30]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][30]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][30]_i_11 
       (.I0(\syncrregs.r[hrdatas][30]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][30]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][30]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][30]_i_12 
       (.I0(\syncrregs.r[hrdatas][30]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][30]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][30]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][30]_i_13 
       (.I0(\syncrregs.r[hrdatas][30]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][30]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][30]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][30]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][30]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][30]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][30]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][30]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][30]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][30]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][30]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][30]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][30]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][30]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][30]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][30]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][30]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][30]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][30]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][30]_i_6 
       (.I0(\syncrregs.r[hrdatas][30]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][30]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][30]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][30]_i_7 
       (.I0(\syncrregs.r[hrdatas][30]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][30]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][30]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][30]_i_8 
       (.I0(\syncrregs.r[hrdatas][30]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][30]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][30]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][30]_i_9 
       (.I0(\syncrregs.r[hrdatas][30]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][30]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][30]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [31]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [31]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][31]_i_10 
       (.I0(\syncrregs.r[hrdatas][31]_i_19_n_0 ),
        .I1(\syncrregs.r[hrdatas][31]_i_20_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][31]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][31]_i_11 
       (.I0(\syncrregs.r[hrdatas][31]_i_21_n_0 ),
        .I1(\syncrregs.r[hrdatas][31]_i_22_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][31]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][31]_i_12 
       (.I0(\syncrregs.r[hrdatas][31]_i_23_n_0 ),
        .I1(\syncrregs.r[hrdatas][31]_i_24_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][31]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][31]_i_13 
       (.I0(\syncrregs.r[hrdatas][31]_i_25_n_0 ),
        .I1(\syncrregs.r[hrdatas][31]_i_26_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][31]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][31]_i_14 
       (.I0(\syncrregs.r[hrdatas][31]_i_27_n_0 ),
        .I1(\syncrregs.r[hrdatas][31]_i_28_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][31]_i_14_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][31]_i_15 
       (.I0(\syncrregs.r[hrdatas][31]_i_29_n_0 ),
        .I1(\syncrregs.r[hrdatas][31]_i_30_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][31]_i_15_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][31]_i_16 
       (.I0(\syncrregs.r[hrdatas][31]_i_31_n_0 ),
        .I1(\syncrregs.r[hrdatas][31]_i_32_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][31]_i_16_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][31]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][31]_i_9_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][31]_i_10_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][31]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][31]_i_6 
       (.I0(\syncrregs.r_reg[hrdatas][31]_i_11_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][31]_i_12_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][31]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][31]_i_7 
       (.I0(\syncrregs.r_reg[hrdatas][31]_i_13_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][31]_i_14_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][31]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][31]_i_8 
       (.I0(\syncrregs.r_reg[hrdatas][31]_i_15_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][31]_i_16_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][31]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][31]_i_9 
       (.I0(\syncrregs.r[hrdatas][31]_i_17_n_0 ),
        .I1(\syncrregs.r[hrdatas][31]_i_18_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][31]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [3]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [3]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][3]_i_10 
       (.I0(\syncrregs.r[hrdatas][3]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][3]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][3]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][3]_i_11 
       (.I0(\syncrregs.r[hrdatas][3]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][3]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][3]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][3]_i_12 
       (.I0(\syncrregs.r[hrdatas][3]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][3]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][3]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][3]_i_13 
       (.I0(\syncrregs.r[hrdatas][3]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][3]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][3]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][3]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][3]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][3]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][3]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][3]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][3]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][3]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][3]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][3]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][3]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][3]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][3]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][3]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][3]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][3]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][3]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][3]_i_6 
       (.I0(\syncrregs.r[hrdatas][3]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][3]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][3]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][3]_i_7 
       (.I0(\syncrregs.r[hrdatas][3]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][3]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][3]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][3]_i_8 
       (.I0(\syncrregs.r[hrdatas][3]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][3]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][3]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][3]_i_9 
       (.I0(\syncrregs.r[hrdatas][3]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][3]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][3]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [4]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [4]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][4]_i_10 
       (.I0(\syncrregs.r[hrdatas][4]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][4]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][4]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][4]_i_11 
       (.I0(\syncrregs.r[hrdatas][4]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][4]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][4]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][4]_i_12 
       (.I0(\syncrregs.r[hrdatas][4]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][4]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][4]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][4]_i_13 
       (.I0(\syncrregs.r[hrdatas][4]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][4]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][4]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][4]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][4]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][4]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][4]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][4]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][4]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][4]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][4]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][4]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][4]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][4]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][4]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][4]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][4]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][4]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][4]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][4]_i_6 
       (.I0(\syncrregs.r[hrdatas][4]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][4]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][4]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][4]_i_7 
       (.I0(\syncrregs.r[hrdatas][4]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][4]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][4]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][4]_i_8 
       (.I0(\syncrregs.r[hrdatas][4]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][4]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][4]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][4]_i_9 
       (.I0(\syncrregs.r[hrdatas][4]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][4]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][4]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r[hrdatas][5]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatas]__0 [5]),
        .S(\v[hrdatas] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][5]_i_10 
       (.I0(\syncrregs.r[hrdatas][5]_i_23_n_0 ),
        .I1(\syncrregs.r[hrdatas][5]_i_24_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][5]_i_10_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][5]_i_11 
       (.I0(\syncrregs.r[hrdatas][5]_i_25_n_0 ),
        .I1(\syncrregs.r[hrdatas][5]_i_26_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][5]_i_11_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][5]_i_12 
       (.I0(\syncrregs.r[hrdatas][5]_i_27_n_0 ),
        .I1(\syncrregs.r[hrdatas][5]_i_28_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][5]_i_12_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][5]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][5]_i_9_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][5]_i_10_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][5]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][5]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][5]_i_11_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][5]_i_12_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][5]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][5]_i_5 
       (.I0(\syncrregs.r[hrdatas][5]_i_13_n_0 ),
        .I1(\syncrregs.r[hrdatas][5]_i_14_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][5]_i_5_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][5]_i_6 
       (.I0(\syncrregs.r[hrdatas][5]_i_15_n_0 ),
        .I1(\syncrregs.r[hrdatas][5]_i_16_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][5]_i_6_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][5]_i_7 
       (.I0(\syncrregs.r[hrdatas][5]_i_17_n_0 ),
        .I1(\syncrregs.r[hrdatas][5]_i_18_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][5]_i_7_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][5]_i_8 
       (.I0(\syncrregs.r[hrdatas][5]_i_19_n_0 ),
        .I1(\syncrregs.r[hrdatas][5]_i_20_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][5]_i_8_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][5]_i_9 
       (.I0(\syncrregs.r[hrdatas][5]_i_21_n_0 ),
        .I1(\syncrregs.r[hrdatas][5]_i_22_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][5]_i_9_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\syncrregs.r[hrdatas][6]_i_1_n_0 ),
        .Q(\syncrregs.r_reg[hrdatas]__0 [6]),
        .S(\v[hrdatas] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][6]_i_10 
       (.I0(\syncrregs.r[hrdatas][6]_i_23_n_0 ),
        .I1(\syncrregs.r[hrdatas][6]_i_24_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][6]_i_10_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][6]_i_11 
       (.I0(\syncrregs.r[hrdatas][6]_i_25_n_0 ),
        .I1(\syncrregs.r[hrdatas][6]_i_26_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][6]_i_11_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][6]_i_12 
       (.I0(\syncrregs.r[hrdatas][6]_i_27_n_0 ),
        .I1(\syncrregs.r[hrdatas][6]_i_28_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][6]_i_12_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][6]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][6]_i_9_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][6]_i_10_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][6]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][6]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][6]_i_11_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][6]_i_12_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][6]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][6]_i_5 
       (.I0(\syncrregs.r[hrdatas][6]_i_13_n_0 ),
        .I1(\syncrregs.r[hrdatas][6]_i_14_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][6]_i_5_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][6]_i_6 
       (.I0(\syncrregs.r[hrdatas][6]_i_15_n_0 ),
        .I1(\syncrregs.r[hrdatas][6]_i_16_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][6]_i_6_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][6]_i_7 
       (.I0(\syncrregs.r[hrdatas][6]_i_17_n_0 ),
        .I1(\syncrregs.r[hrdatas][6]_i_18_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][6]_i_7_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][6]_i_8 
       (.I0(\syncrregs.r[hrdatas][6]_i_19_n_0 ),
        .I1(\syncrregs.r[hrdatas][6]_i_20_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][6]_i_8_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][6]_i_9 
       (.I0(\syncrregs.r[hrdatas][6]_i_21_n_0 ),
        .I1(\syncrregs.r[hrdatas][6]_i_22_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][6]_i_9_n_0 ),
        .S(sel0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [7]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [7]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][7]_i_10 
       (.I0(\syncrregs.r[hrdatas][7]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][7]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][7]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][7]_i_11 
       (.I0(\syncrregs.r[hrdatas][7]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][7]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][7]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][7]_i_12 
       (.I0(\syncrregs.r[hrdatas][7]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][7]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][7]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][7]_i_13 
       (.I0(\syncrregs.r[hrdatas][7]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][7]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][7]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][7]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][7]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][7]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][7]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][7]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][7]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][7]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][7]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][7]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][7]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][7]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][7]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][7]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][7]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][7]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][7]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][7]_i_6 
       (.I0(\syncrregs.r[hrdatas][7]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][7]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][7]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][7]_i_7 
       (.I0(\syncrregs.r[hrdatas][7]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][7]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][7]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][7]_i_8 
       (.I0(\syncrregs.r[hrdatas][7]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][7]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][7]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][7]_i_9 
       (.I0(\syncrregs.r[hrdatas][7]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][7]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][7]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [8]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [8]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][8]_i_10 
       (.I0(\syncrregs.r[hrdatas][8]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][8]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][8]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][8]_i_11 
       (.I0(\syncrregs.r[hrdatas][8]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][8]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][8]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][8]_i_12 
       (.I0(\syncrregs.r[hrdatas][8]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][8]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][8]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][8]_i_13 
       (.I0(\syncrregs.r[hrdatas][8]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][8]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][8]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][8]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][8]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][8]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][8]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][8]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][8]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][8]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][8]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][8]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][8]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][8]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][8]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][8]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][8]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][8]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][8]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][8]_i_6 
       (.I0(\syncrregs.r[hrdatas][8]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][8]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][8]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][8]_i_7 
       (.I0(\syncrregs.r[hrdatas][8]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][8]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][8]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][8]_i_8 
       (.I0(\syncrregs.r[hrdatas][8]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][8]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][8]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][8]_i_9 
       (.I0(\syncrregs.r[hrdatas][8]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][8]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][8]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hrdatas][9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\slvo[15][hready]__0 [9]),
        .Q(\syncrregs.r_reg[hrdatas]__0 [9]),
        .R(\v[hrdatas] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][9]_i_10 
       (.I0(\syncrregs.r[hrdatas][9]_i_22_n_0 ),
        .I1(\syncrregs.r[hrdatas][9]_i_23_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][9]_i_10_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][9]_i_11 
       (.I0(\syncrregs.r[hrdatas][9]_i_24_n_0 ),
        .I1(\syncrregs.r[hrdatas][9]_i_25_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][9]_i_11_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][9]_i_12 
       (.I0(\syncrregs.r[hrdatas][9]_i_26_n_0 ),
        .I1(\syncrregs.r[hrdatas][9]_i_27_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][9]_i_12_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][9]_i_13 
       (.I0(\syncrregs.r[hrdatas][9]_i_28_n_0 ),
        .I1(\syncrregs.r[hrdatas][9]_i_29_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][9]_i_13_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][9]_i_2 
       (.I0(\syncrregs.r_reg[hrdatas][9]_i_6_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][9]_i_7_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][9]_i_2_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][9]_i_3 
       (.I0(\syncrregs.r_reg[hrdatas][9]_i_8_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][9]_i_9_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][9]_i_3_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][9]_i_4 
       (.I0(\syncrregs.r_reg[hrdatas][9]_i_10_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][9]_i_11_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][9]_i_4_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \syncrregs.r_reg[hrdatas][9]_i_5 
       (.I0(\syncrregs.r_reg[hrdatas][9]_i_12_n_0 ),
        .I1(\syncrregs.r_reg[hrdatas][9]_i_13_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][9]_i_5_n_0 ),
        .S(\syncrregs.r_reg[haddr_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][9]_i_6 
       (.I0(\syncrregs.r[hrdatas][9]_i_14_n_0 ),
        .I1(\syncrregs.r[hrdatas][9]_i_15_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][9]_i_6_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][9]_i_7 
       (.I0(\syncrregs.r[hrdatas][9]_i_16_n_0 ),
        .I1(\syncrregs.r[hrdatas][9]_i_17_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][9]_i_7_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][9]_i_8 
       (.I0(\syncrregs.r[hrdatas][9]_i_18_n_0 ),
        .I1(\syncrregs.r[hrdatas][9]_i_19_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][9]_i_8_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \syncrregs.r_reg[hrdatas][9]_i_9 
       (.I0(\syncrregs.r[hrdatas][9]_i_20_n_0 ),
        .I1(\syncrregs.r[hrdatas][9]_i_21_n_0 ),
        .O(\syncrregs.r_reg[hrdatas][9]_i_9_n_0 ),
        .S(\syncrregs.r_reg[haddr][7]_rep_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hready] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(rin),
        .Q(\syncrregs.r_reg[hready_n_0_] ),
        .R(slvi));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hslave][0] 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(p_6_out),
        .Q(\syncrregs.r_reg[hslave]__0 [0]),
        .R(\syncrregs.r[htrans][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hslave][1] 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(p_11_out),
        .Q(\syncrregs.r_reg[hslave]__0 [1]),
        .R(\syncrregs.r[htrans][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[hslave][2] 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(p_14_out),
        .Q(\syncrregs.r_reg[hslave]__0 [2]),
        .R(\syncrregs.r[htrans][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \syncrregs.r_reg[htrans][1] 
       (.C(clk),
        .CE(\slvi[hready] ),
        .D(\slvi[htrans] [1]),
        .Q(\syncrregs.r_reg[htrans_n_0_][1] ),
        .R(\syncrregs.r[htrans][1]_i_1_n_0 ));
endmodule
