module tiny_encryption_algorithm
   (clock,
    reset,
    start,
    ready,
    key,
    text,
    backdoor,
    cipher);
  output backdoor;
  input clock;
  input reset;
  input start;
  output ready;
  input [127:0]key;
  input [63:0]text;
  output [63:0]cipher;

  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const0>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const1>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:0]cipher;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire clock;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cnt;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cnt[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cnt[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cnt[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cnt[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cnt[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cnt[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cnt[6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cnt[6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cnt_reg_n_0_;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cnt_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cnt_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cnt_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cnt_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire feistelKey0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]feistelKey0__0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:27]feistelKey1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]k0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]k1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]k2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]k3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]key;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]p_0_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]plusOp;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:3]plusOp0_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]plusOp1_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ready;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire reset;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sel;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire start;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sum;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum[12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum[12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum[12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum[16]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum[16]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum[16]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum[20]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum[20]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum[24]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum[24]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum[24]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum[28]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum[28]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum[4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum[4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum[8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]sum_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[0]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[0]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[0]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[0]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[0]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[0]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[0]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[12]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[12]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[12]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[12]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[12]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[12]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[12]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[16]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[16]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[16]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[16]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[16]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[16]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[16]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[20]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[20]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[20]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[20]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[20]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[20]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[20]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[24]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[24]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[24]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[24]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[24]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[24]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[24]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[28]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[28]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[28]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[28]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[4]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[4]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[4]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[4]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[4]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[4]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[4]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[8]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[8]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[8]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[8]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[8]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[8]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sum_reg[8]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:0]text;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire v1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[11]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[11]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[11]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[11]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[11]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[11]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[11]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[11]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[11]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[11]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[11]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[11]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[11]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[11]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[11]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[11]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[15]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[15]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[15]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[15]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[15]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[15]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[15]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[15]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[15]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[15]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[15]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[15]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[15]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[15]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[15]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[15]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[15]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[19]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[19]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[19]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[19]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[19]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[19]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[19]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[19]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[19]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[19]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[19]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[19]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[19]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[19]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[19]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[19]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[19]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[19]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[19]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[19]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[23]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[23]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[23]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[23]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[23]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[23]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[23]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[23]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[23]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[23]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[23]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[23]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[23]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[23]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[23]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[23]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[23]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[23]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[23]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[23]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[27]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[27]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[27]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[27]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[27]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[27]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[27]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[27]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[27]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[27]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[27]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[27]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[27]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[27]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[27]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[27]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[27]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[27]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[27]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[31]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[31]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[31]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[31]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[31]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[31]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[31]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[31]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[31]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[31]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[31]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[31]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[31]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[3]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[3]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[3]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[3]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[3]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[3]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[3]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[3]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[7]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[7]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[7]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[7]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[7]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[7]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[7]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[7]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[7]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[7]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[7]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[7]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[7]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[7]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[7]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1[7]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]v1_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[11]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[11]_i_11_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[11]_i_11_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[11]_i_11_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[11]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[11]_i_12_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[11]_i_12_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[11]_i_12_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[11]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[11]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[11]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[11]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[11]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[11]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[11]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[15]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[15]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[15]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[15]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[15]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[15]_i_11_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[15]_i_11_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[15]_i_11_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[15]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[15]_i_12_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[15]_i_12_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[15]_i_12_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[15]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[15]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[15]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[15]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[15]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[15]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[15]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[19]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[19]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[19]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[19]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[19]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[19]_i_11_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[19]_i_11_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[19]_i_11_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[19]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[19]_i_12_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[19]_i_12_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[19]_i_12_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[19]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[19]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[19]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[19]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[19]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[19]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[19]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[23]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[23]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[23]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[23]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[23]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[23]_i_11_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[23]_i_11_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[23]_i_11_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[23]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[23]_i_12_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[23]_i_12_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[23]_i_12_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[23]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[23]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[23]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[23]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[23]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[23]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[23]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[27]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[27]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[27]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[27]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[27]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[27]_i_11_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[27]_i_11_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[27]_i_11_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[27]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[27]_i_12_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[27]_i_12_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[27]_i_12_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[27]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[27]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[27]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[27]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[27]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[27]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[27]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[31]_i_12_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[31]_i_12_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[31]_i_12_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[31]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[31]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[31]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[31]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[31]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[31]_i_9_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[31]_i_9_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[31]_i_9_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[3]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[3]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[3]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[3]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[3]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[3]_i_11_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[3]_i_11_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[3]_i_11_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[3]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[3]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[3]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[3]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[3]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[3]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[3]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[7]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[7]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[7]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[7]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[7]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[7]_i_11_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[7]_i_11_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[7]_i_11_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[7]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[7]_i_12_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[7]_i_12_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[7]_i_12_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[7]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[7]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[7]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[7]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[7]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[7]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v1_reg[7]_i_1_n_7 ;

  assign backdoor =  v1 ;

  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND
       (.G(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC
       (.P(\<const1>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cnt[0]_i_1 
       (.I0(sel),
        .I1(ready),
        .O(cnt));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \cnt[1]_i_1 
       (.I0(cnt_reg_n_0_),
        .I1(sel),
        .I2(ready),
        .O(\cnt[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair0" *) 
  LUT4 #(
    .INIT(16'h006A)) 
    \cnt[2]_i_1 
       (.I0(\cnt_reg_n_0_[2] ),
        .I1(cnt_reg_n_0_),
        .I2(sel),
        .I3(ready),
        .O(\cnt[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair0" *) 
  LUT5 #(
    .INIT(32'h00006AAA)) 
    \cnt[3]_i_1 
       (.I0(\cnt_reg_n_0_[3] ),
        .I1(\cnt_reg_n_0_[2] ),
        .I2(sel),
        .I3(cnt_reg_n_0_),
        .I4(ready),
        .O(\cnt[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000006AAAAAAA)) 
    \cnt[4]_i_1 
       (.I0(\cnt_reg_n_0_[4] ),
        .I1(\cnt_reg_n_0_[3] ),
        .I2(cnt_reg_n_0_),
        .I3(sel),
        .I4(\cnt_reg_n_0_[2] ),
        .I5(ready),
        .O(\cnt[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair19" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \cnt[5]_i_1 
       (.I0(\cnt_reg_n_0_[5] ),
        .I1(\cnt[6]_i_3_n_0 ),
        .I2(ready),
        .O(\cnt[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \cnt[6]_i_1 
       (.I0(start),
        .I1(ready),
        .O(\cnt[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair19" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \cnt[6]_i_2 
       (.I0(\cnt_reg_n_0_[5] ),
        .I1(\cnt[6]_i_3_n_0 ),
        .I2(ready),
        .O(\cnt[6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h80000000)) 
    \cnt[6]_i_3 
       (.I0(\cnt_reg_n_0_[4] ),
        .I1(\cnt_reg_n_0_[2] ),
        .I2(sel),
        .I3(cnt_reg_n_0_),
        .I4(\cnt_reg_n_0_[3] ),
        .O(\cnt[6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \cnt_reg[0] 
       (.C(clock),
        .CE(\cnt[6]_i_1_n_0 ),
        .D(cnt),
        .Q(sel),
        .S(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \cnt_reg[1] 
       (.C(clock),
        .CE(\cnt[6]_i_1_n_0 ),
        .D(\cnt[1]_i_1_n_0 ),
        .Q(cnt_reg_n_0_),
        .S(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \cnt_reg[2] 
       (.C(clock),
        .CE(\cnt[6]_i_1_n_0 ),
        .D(\cnt[2]_i_1_n_0 ),
        .Q(\cnt_reg_n_0_[2] ),
        .S(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \cnt_reg[3] 
       (.C(clock),
        .CE(\cnt[6]_i_1_n_0 ),
        .D(\cnt[3]_i_1_n_0 ),
        .Q(\cnt_reg_n_0_[3] ),
        .S(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \cnt_reg[4] 
       (.C(clock),
        .CE(\cnt[6]_i_1_n_0 ),
        .D(\cnt[4]_i_1_n_0 ),
        .Q(\cnt_reg_n_0_[4] ),
        .S(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \cnt_reg[5] 
       (.C(clock),
        .CE(\cnt[6]_i_1_n_0 ),
        .D(\cnt[5]_i_1_n_0 ),
        .Q(\cnt_reg_n_0_[5] ),
        .S(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \cnt_reg[6] 
       (.C(clock),
        .CE(\cnt[6]_i_1_n_0 ),
        .D(\cnt[6]_i_2_n_0 ),
        .Q(ready),
        .S(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[0] 
       (.C(clock),
        .CE(ready),
        .D(key[0]),
        .Q(k0[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[10] 
       (.C(clock),
        .CE(ready),
        .D(key[10]),
        .Q(k0[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[11] 
       (.C(clock),
        .CE(ready),
        .D(key[11]),
        .Q(k0[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[12] 
       (.C(clock),
        .CE(ready),
        .D(key[12]),
        .Q(k0[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[13] 
       (.C(clock),
        .CE(ready),
        .D(key[13]),
        .Q(k0[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[14] 
       (.C(clock),
        .CE(ready),
        .D(key[14]),
        .Q(k0[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[15] 
       (.C(clock),
        .CE(ready),
        .D(key[15]),
        .Q(k0[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[16] 
       (.C(clock),
        .CE(ready),
        .D(key[16]),
        .Q(k0[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[17] 
       (.C(clock),
        .CE(ready),
        .D(key[17]),
        .Q(k0[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[18] 
       (.C(clock),
        .CE(ready),
        .D(key[18]),
        .Q(k0[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[19] 
       (.C(clock),
        .CE(ready),
        .D(key[19]),
        .Q(k0[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[1] 
       (.C(clock),
        .CE(ready),
        .D(key[1]),
        .Q(k0[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[20] 
       (.C(clock),
        .CE(ready),
        .D(key[20]),
        .Q(k0[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[21] 
       (.C(clock),
        .CE(ready),
        .D(key[21]),
        .Q(k0[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[22] 
       (.C(clock),
        .CE(ready),
        .D(key[22]),
        .Q(k0[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[23] 
       (.C(clock),
        .CE(ready),
        .D(key[23]),
        .Q(k0[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[24] 
       (.C(clock),
        .CE(ready),
        .D(key[24]),
        .Q(k0[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[25] 
       (.C(clock),
        .CE(ready),
        .D(key[25]),
        .Q(k0[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[26] 
       (.C(clock),
        .CE(ready),
        .D(key[26]),
        .Q(k0[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[27] 
       (.C(clock),
        .CE(ready),
        .D(key[27]),
        .Q(k0[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[28] 
       (.C(clock),
        .CE(ready),
        .D(key[28]),
        .Q(k0[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[29] 
       (.C(clock),
        .CE(ready),
        .D(key[29]),
        .Q(k0[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[2] 
       (.C(clock),
        .CE(ready),
        .D(key[2]),
        .Q(k0[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[30] 
       (.C(clock),
        .CE(ready),
        .D(key[30]),
        .Q(k0[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[31] 
       (.C(clock),
        .CE(ready),
        .D(key[31]),
        .Q(k0[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[3] 
       (.C(clock),
        .CE(ready),
        .D(key[3]),
        .Q(k0[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[4] 
       (.C(clock),
        .CE(ready),
        .D(key[4]),
        .Q(k0[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[5] 
       (.C(clock),
        .CE(ready),
        .D(key[5]),
        .Q(k0[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[6] 
       (.C(clock),
        .CE(ready),
        .D(key[6]),
        .Q(k0[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[7] 
       (.C(clock),
        .CE(ready),
        .D(key[7]),
        .Q(k0[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[8] 
       (.C(clock),
        .CE(ready),
        .D(key[8]),
        .Q(k0[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[9] 
       (.C(clock),
        .CE(ready),
        .D(key[9]),
        .Q(k0[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[0] 
       (.C(clock),
        .CE(ready),
        .D(key[32]),
        .Q(k1[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[10] 
       (.C(clock),
        .CE(ready),
        .D(key[42]),
        .Q(k1[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[11] 
       (.C(clock),
        .CE(ready),
        .D(key[43]),
        .Q(k1[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[12] 
       (.C(clock),
        .CE(ready),
        .D(key[44]),
        .Q(k1[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[13] 
       (.C(clock),
        .CE(ready),
        .D(key[45]),
        .Q(k1[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[14] 
       (.C(clock),
        .CE(ready),
        .D(key[46]),
        .Q(k1[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[15] 
       (.C(clock),
        .CE(ready),
        .D(key[47]),
        .Q(k1[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[16] 
       (.C(clock),
        .CE(ready),
        .D(key[48]),
        .Q(k1[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[17] 
       (.C(clock),
        .CE(ready),
        .D(key[49]),
        .Q(k1[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[18] 
       (.C(clock),
        .CE(ready),
        .D(key[50]),
        .Q(k1[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[19] 
       (.C(clock),
        .CE(ready),
        .D(key[51]),
        .Q(k1[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[1] 
       (.C(clock),
        .CE(ready),
        .D(key[33]),
        .Q(k1[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[20] 
       (.C(clock),
        .CE(ready),
        .D(key[52]),
        .Q(k1[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[21] 
       (.C(clock),
        .CE(ready),
        .D(key[53]),
        .Q(k1[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[22] 
       (.C(clock),
        .CE(ready),
        .D(key[54]),
        .Q(k1[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[23] 
       (.C(clock),
        .CE(ready),
        .D(key[55]),
        .Q(k1[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[24] 
       (.C(clock),
        .CE(ready),
        .D(key[56]),
        .Q(k1[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[25] 
       (.C(clock),
        .CE(ready),
        .D(key[57]),
        .Q(k1[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[26] 
       (.C(clock),
        .CE(ready),
        .D(key[58]),
        .Q(k1[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[27] 
       (.C(clock),
        .CE(ready),
        .D(key[59]),
        .Q(k1[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[28] 
       (.C(clock),
        .CE(ready),
        .D(key[60]),
        .Q(k1[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[29] 
       (.C(clock),
        .CE(ready),
        .D(key[61]),
        .Q(k1[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[2] 
       (.C(clock),
        .CE(ready),
        .D(key[34]),
        .Q(k1[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[30] 
       (.C(clock),
        .CE(ready),
        .D(key[62]),
        .Q(k1[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[31] 
       (.C(clock),
        .CE(ready),
        .D(key[63]),
        .Q(k1[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[3] 
       (.C(clock),
        .CE(ready),
        .D(key[35]),
        .Q(k1[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[4] 
       (.C(clock),
        .CE(ready),
        .D(key[36]),
        .Q(k1[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[5] 
       (.C(clock),
        .CE(ready),
        .D(key[37]),
        .Q(k1[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[6] 
       (.C(clock),
        .CE(ready),
        .D(key[38]),
        .Q(k1[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[7] 
       (.C(clock),
        .CE(ready),
        .D(key[39]),
        .Q(k1[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[8] 
       (.C(clock),
        .CE(ready),
        .D(key[40]),
        .Q(k1[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k1_reg[9] 
       (.C(clock),
        .CE(ready),
        .D(key[41]),
        .Q(k1[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[0] 
       (.C(clock),
        .CE(ready),
        .D(key[64]),
        .Q(k2[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[10] 
       (.C(clock),
        .CE(ready),
        .D(key[74]),
        .Q(k2[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[11] 
       (.C(clock),
        .CE(ready),
        .D(key[75]),
        .Q(k2[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[12] 
       (.C(clock),
        .CE(ready),
        .D(key[76]),
        .Q(k2[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[13] 
       (.C(clock),
        .CE(ready),
        .D(key[77]),
        .Q(k2[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[14] 
       (.C(clock),
        .CE(ready),
        .D(key[78]),
        .Q(k2[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[15] 
       (.C(clock),
        .CE(ready),
        .D(key[79]),
        .Q(k2[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[16] 
       (.C(clock),
        .CE(ready),
        .D(key[80]),
        .Q(k2[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[17] 
       (.C(clock),
        .CE(ready),
        .D(key[81]),
        .Q(k2[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[18] 
       (.C(clock),
        .CE(ready),
        .D(key[82]),
        .Q(k2[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[19] 
       (.C(clock),
        .CE(ready),
        .D(key[83]),
        .Q(k2[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[1] 
       (.C(clock),
        .CE(ready),
        .D(key[65]),
        .Q(k2[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[20] 
       (.C(clock),
        .CE(ready),
        .D(key[84]),
        .Q(k2[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[21] 
       (.C(clock),
        .CE(ready),
        .D(key[85]),
        .Q(k2[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[22] 
       (.C(clock),
        .CE(ready),
        .D(key[86]),
        .Q(k2[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[23] 
       (.C(clock),
        .CE(ready),
        .D(key[87]),
        .Q(k2[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[24] 
       (.C(clock),
        .CE(ready),
        .D(key[88]),
        .Q(k2[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[25] 
       (.C(clock),
        .CE(ready),
        .D(key[89]),
        .Q(k2[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[26] 
       (.C(clock),
        .CE(ready),
        .D(key[90]),
        .Q(k2[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[27] 
       (.C(clock),
        .CE(ready),
        .D(key[91]),
        .Q(k2[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[28] 
       (.C(clock),
        .CE(ready),
        .D(key[92]),
        .Q(k2[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[29] 
       (.C(clock),
        .CE(ready),
        .D(key[93]),
        .Q(k2[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[2] 
       (.C(clock),
        .CE(ready),
        .D(key[66]),
        .Q(k2[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[30] 
       (.C(clock),
        .CE(ready),
        .D(key[94]),
        .Q(k2[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[31] 
       (.C(clock),
        .CE(ready),
        .D(key[95]),
        .Q(k2[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[3] 
       (.C(clock),
        .CE(ready),
        .D(key[67]),
        .Q(k2[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[4] 
       (.C(clock),
        .CE(ready),
        .D(key[68]),
        .Q(k2[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[5] 
       (.C(clock),
        .CE(ready),
        .D(key[69]),
        .Q(k2[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[6] 
       (.C(clock),
        .CE(ready),
        .D(key[70]),
        .Q(k2[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[7] 
       (.C(clock),
        .CE(ready),
        .D(key[71]),
        .Q(k2[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[8] 
       (.C(clock),
        .CE(ready),
        .D(key[72]),
        .Q(k2[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k2_reg[9] 
       (.C(clock),
        .CE(ready),
        .D(key[73]),
        .Q(k2[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[0] 
       (.C(clock),
        .CE(ready),
        .D(key[96]),
        .Q(k3[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[10] 
       (.C(clock),
        .CE(ready),
        .D(key[106]),
        .Q(k3[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[11] 
       (.C(clock),
        .CE(ready),
        .D(key[107]),
        .Q(k3[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[12] 
       (.C(clock),
        .CE(ready),
        .D(key[108]),
        .Q(k3[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[13] 
       (.C(clock),
        .CE(ready),
        .D(key[109]),
        .Q(k3[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[14] 
       (.C(clock),
        .CE(ready),
        .D(key[110]),
        .Q(k3[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[15] 
       (.C(clock),
        .CE(ready),
        .D(key[111]),
        .Q(k3[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[16] 
       (.C(clock),
        .CE(ready),
        .D(key[112]),
        .Q(k3[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[17] 
       (.C(clock),
        .CE(ready),
        .D(key[113]),
        .Q(k3[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[18] 
       (.C(clock),
        .CE(ready),
        .D(key[114]),
        .Q(k3[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[19] 
       (.C(clock),
        .CE(ready),
        .D(key[115]),
        .Q(k3[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[1] 
       (.C(clock),
        .CE(ready),
        .D(key[97]),
        .Q(k3[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[20] 
       (.C(clock),
        .CE(ready),
        .D(key[116]),
        .Q(k3[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[21] 
       (.C(clock),
        .CE(ready),
        .D(key[117]),
        .Q(k3[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[22] 
       (.C(clock),
        .CE(ready),
        .D(key[118]),
        .Q(k3[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[23] 
       (.C(clock),
        .CE(ready),
        .D(key[119]),
        .Q(k3[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[24] 
       (.C(clock),
        .CE(ready),
        .D(key[120]),
        .Q(k3[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[25] 
       (.C(clock),
        .CE(ready),
        .D(key[121]),
        .Q(k3[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[26] 
       (.C(clock),
        .CE(ready),
        .D(key[122]),
        .Q(k3[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[27] 
       (.C(clock),
        .CE(ready),
        .D(key[123]),
        .Q(k3[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[28] 
       (.C(clock),
        .CE(ready),
        .D(key[124]),
        .Q(k3[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[29] 
       (.C(clock),
        .CE(ready),
        .D(key[125]),
        .Q(k3[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[2] 
       (.C(clock),
        .CE(ready),
        .D(key[98]),
        .Q(k3[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[30] 
       (.C(clock),
        .CE(ready),
        .D(key[126]),
        .Q(k3[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[31] 
       (.C(clock),
        .CE(ready),
        .D(key[127]),
        .Q(k3[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[3] 
       (.C(clock),
        .CE(ready),
        .D(key[99]),
        .Q(k3[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[4] 
       (.C(clock),
        .CE(ready),
        .D(key[100]),
        .Q(k3[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[5] 
       (.C(clock),
        .CE(ready),
        .D(key[101]),
        .Q(k3[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[6] 
       (.C(clock),
        .CE(ready),
        .D(key[102]),
        .Q(k3[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[7] 
       (.C(clock),
        .CE(ready),
        .D(key[103]),
        .Q(k3[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[8] 
       (.C(clock),
        .CE(ready),
        .D(key[104]),
        .Q(k3[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k3_reg[9] 
       (.C(clock),
        .CE(ready),
        .D(key[105]),
        .Q(k3[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \sum[0]_i_2 
       (.I0(sum_reg[3]),
        .O(sum));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \sum[0]_i_5 
       (.I0(sum_reg[0]),
        .O(\sum[0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \sum[12]_i_3 
       (.I0(sum_reg[14]),
        .O(\sum[12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \sum[12]_i_4 
       (.I0(sum_reg[13]),
        .O(\sum[12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \sum[12]_i_5 
       (.I0(sum_reg[12]),
        .O(\sum[12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \sum[16]_i_3 
       (.I0(sum_reg[18]),
        .O(\sum[16]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \sum[16]_i_4 
       (.I0(sum_reg[17]),
        .O(\sum[16]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \sum[16]_i_5 
       (.I0(sum_reg[16]),
        .O(\sum[16]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \sum[20]_i_4 
       (.I0(sum_reg[21]),
        .O(\sum[20]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \sum[20]_i_5 
       (.I0(sum_reg[20]),
        .O(\sum[20]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \sum[24]_i_2 
       (.I0(sum_reg[27]),
        .O(\sum[24]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \sum[24]_i_3 
       (.I0(sum_reg[26]),
        .O(\sum[24]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \sum[24]_i_4 
       (.I0(sum_reg[25]),
        .O(\sum[24]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \sum[28]_i_2 
       (.I0(sum_reg[31]),
        .O(\sum[28]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \sum[28]_i_5 
       (.I0(sum_reg[28]),
        .O(\sum[28]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \sum[4]_i_2 
       (.I0(sum_reg[7]),
        .O(\sum[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \sum[4]_i_4 
       (.I0(sum_reg[5]),
        .O(\sum[4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \sum[4]_i_5 
       (.I0(sum_reg[4]),
        .O(\sum[4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \sum[8]_i_2 
       (.I0(sum_reg[11]),
        .O(\sum[8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \sum[8]_i_5 
       (.I0(sum_reg[8]),
        .O(\sum[8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \sum_reg[0] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[0]_i_1_n_7 ),
        .Q(sum_reg[0]),
        .S(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \sum_reg[0]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO({\sum_reg[0]_i_1_n_0 ,\sum_reg[0]_i_1_n_1 ,\sum_reg[0]_i_1_n_2 ,\sum_reg[0]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .O({\sum_reg[0]_i_1_n_4 ,\sum_reg[0]_i_1_n_5 ,\sum_reg[0]_i_1_n_6 ,\sum_reg[0]_i_1_n_7 }),
        .S({sum,sum_reg[2:1],\sum[0]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \sum_reg[10] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[8]_i_1_n_5 ),
        .Q(sum_reg[10]),
        .R(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \sum_reg[11] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[8]_i_1_n_4 ),
        .Q(sum_reg[11]),
        .S(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \sum_reg[12] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[12]_i_1_n_7 ),
        .Q(sum_reg[12]),
        .S(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \sum_reg[12]_i_1 
       (.CI(\sum_reg[8]_i_1_n_0 ),
        .CO({\sum_reg[12]_i_1_n_0 ,\sum_reg[12]_i_1_n_1 ,\sum_reg[12]_i_1_n_2 ,\sum_reg[12]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .O({\sum_reg[12]_i_1_n_4 ,\sum_reg[12]_i_1_n_5 ,\sum_reg[12]_i_1_n_6 ,\sum_reg[12]_i_1_n_7 }),
        .S({sum_reg[15],\sum[12]_i_3_n_0 ,\sum[12]_i_4_n_0 ,\sum[12]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \sum_reg[13] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[12]_i_1_n_6 ),
        .Q(sum_reg[13]),
        .S(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \sum_reg[14] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[12]_i_1_n_5 ),
        .Q(sum_reg[14]),
        .S(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \sum_reg[15] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[12]_i_1_n_4 ),
        .Q(sum_reg[15]),
        .R(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \sum_reg[16] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[16]_i_1_n_7 ),
        .Q(sum_reg[16]),
        .S(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \sum_reg[16]_i_1 
       (.CI(\sum_reg[12]_i_1_n_0 ),
        .CO({\sum_reg[16]_i_1_n_0 ,\sum_reg[16]_i_1_n_1 ,\sum_reg[16]_i_1_n_2 ,\sum_reg[16]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .O({\sum_reg[16]_i_1_n_4 ,\sum_reg[16]_i_1_n_5 ,\sum_reg[16]_i_1_n_6 ,\sum_reg[16]_i_1_n_7 }),
        .S({sum_reg[19],\sum[16]_i_3_n_0 ,\sum[16]_i_4_n_0 ,\sum[16]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \sum_reg[17] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[16]_i_1_n_6 ),
        .Q(sum_reg[17]),
        .S(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \sum_reg[18] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[16]_i_1_n_5 ),
        .Q(sum_reg[18]),
        .S(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \sum_reg[19] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[16]_i_1_n_4 ),
        .Q(sum_reg[19]),
        .R(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \sum_reg[1] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[0]_i_1_n_6 ),
        .Q(sum_reg[1]),
        .R(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \sum_reg[20] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[20]_i_1_n_7 ),
        .Q(sum_reg[20]),
        .S(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \sum_reg[20]_i_1 
       (.CI(\sum_reg[16]_i_1_n_0 ),
        .CO({\sum_reg[20]_i_1_n_0 ,\sum_reg[20]_i_1_n_1 ,\sum_reg[20]_i_1_n_2 ,\sum_reg[20]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .O({\sum_reg[20]_i_1_n_4 ,\sum_reg[20]_i_1_n_5 ,\sum_reg[20]_i_1_n_6 ,\sum_reg[20]_i_1_n_7 }),
        .S({sum_reg[23:22],\sum[20]_i_4_n_0 ,\sum[20]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \sum_reg[21] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[20]_i_1_n_6 ),
        .Q(sum_reg[21]),
        .S(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \sum_reg[22] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[20]_i_1_n_5 ),
        .Q(sum_reg[22]),
        .R(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \sum_reg[23] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[20]_i_1_n_4 ),
        .Q(sum_reg[23]),
        .R(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \sum_reg[24] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[24]_i_1_n_7 ),
        .Q(sum_reg[24]),
        .R(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \sum_reg[24]_i_1 
       (.CI(\sum_reg[20]_i_1_n_0 ),
        .CO({\sum_reg[24]_i_1_n_0 ,\sum_reg[24]_i_1_n_1 ,\sum_reg[24]_i_1_n_2 ,\sum_reg[24]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 }),
        .O({\sum_reg[24]_i_1_n_4 ,\sum_reg[24]_i_1_n_5 ,\sum_reg[24]_i_1_n_6 ,\sum_reg[24]_i_1_n_7 }),
        .S({\sum[24]_i_2_n_0 ,\sum[24]_i_3_n_0 ,\sum[24]_i_4_n_0 ,sum_reg[24]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \sum_reg[25] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[24]_i_1_n_6 ),
        .Q(sum_reg[25]),
        .S(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \sum_reg[26] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[24]_i_1_n_5 ),
        .Q(sum_reg[26]),
        .S(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \sum_reg[27] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[24]_i_1_n_4 ),
        .Q(sum_reg[27]),
        .S(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \sum_reg[28] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[28]_i_1_n_7 ),
        .Q(sum_reg[28]),
        .S(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \sum_reg[28]_i_1 
       (.CI(\sum_reg[24]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .O({\sum_reg[28]_i_1_n_4 ,\sum_reg[28]_i_1_n_5 ,\sum_reg[28]_i_1_n_6 ,\sum_reg[28]_i_1_n_7 }),
        .S({\sum[28]_i_2_n_0 ,sum_reg[30:29],\sum[28]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \sum_reg[29] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[28]_i_1_n_6 ),
        .Q(sum_reg[29]),
        .R(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \sum_reg[2] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[0]_i_1_n_5 ),
        .Q(sum_reg[2]),
        .R(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \sum_reg[30] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[28]_i_1_n_5 ),
        .Q(sum_reg[30]),
        .R(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \sum_reg[31] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[28]_i_1_n_4 ),
        .Q(sum_reg[31]),
        .S(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \sum_reg[3] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[0]_i_1_n_4 ),
        .Q(sum_reg[3]),
        .S(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \sum_reg[4] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[4]_i_1_n_7 ),
        .Q(sum_reg[4]),
        .S(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \sum_reg[4]_i_1 
       (.CI(\sum_reg[0]_i_1_n_0 ),
        .CO({\sum_reg[4]_i_1_n_0 ,\sum_reg[4]_i_1_n_1 ,\sum_reg[4]_i_1_n_2 ,\sum_reg[4]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .O({\sum_reg[4]_i_1_n_4 ,\sum_reg[4]_i_1_n_5 ,\sum_reg[4]_i_1_n_6 ,\sum_reg[4]_i_1_n_7 }),
        .S({\sum[4]_i_2_n_0 ,sum_reg[6],\sum[4]_i_4_n_0 ,\sum[4]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \sum_reg[5] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[4]_i_1_n_6 ),
        .Q(sum_reg[5]),
        .S(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \sum_reg[6] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[4]_i_1_n_5 ),
        .Q(sum_reg[6]),
        .R(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \sum_reg[7] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[4]_i_1_n_4 ),
        .Q(sum_reg[7]),
        .S(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \sum_reg[8] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[8]_i_1_n_7 ),
        .Q(sum_reg[8]),
        .S(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \sum_reg[8]_i_1 
       (.CI(\sum_reg[4]_i_1_n_0 ),
        .CO({\sum_reg[8]_i_1_n_0 ,\sum_reg[8]_i_1_n_1 ,\sum_reg[8]_i_1_n_2 ,\sum_reg[8]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .O({\sum_reg[8]_i_1_n_4 ,\sum_reg[8]_i_1_n_5 ,\sum_reg[8]_i_1_n_6 ,\sum_reg[8]_i_1_n_7 }),
        .S({\sum[8]_i_2_n_0 ,sum_reg[10:9],\sum[8]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \sum_reg[9] 
       (.C(clock),
        .CE(sel),
        .D(\sum_reg[8]_i_1_n_6 ),
        .Q(sum_reg[9]),
        .R(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair1" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[0]_i_1 
       (.I0(text[0]),
        .I1(cipher[32]),
        .I2(ready),
        .O(p_0_in[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[10]_i_1 
       (.I0(text[10]),
        .I1(cipher[42]),
        .I2(ready),
        .O(p_0_in[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[11]_i_1 
       (.I0(text[11]),
        .I1(cipher[43]),
        .I2(ready),
        .O(p_0_in[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[12]_i_1 
       (.I0(text[12]),
        .I1(cipher[44]),
        .I2(ready),
        .O(p_0_in[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[13]_i_1 
       (.I0(text[13]),
        .I1(cipher[45]),
        .I2(ready),
        .O(p_0_in[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[14]_i_1 
       (.I0(text[14]),
        .I1(cipher[46]),
        .I2(ready),
        .O(p_0_in[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[15]_i_1 
       (.I0(text[15]),
        .I1(cipher[47]),
        .I2(ready),
        .O(p_0_in[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair11" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[16]_i_1 
       (.I0(text[16]),
        .I1(cipher[48]),
        .I2(ready),
        .O(p_0_in[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair12" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[17]_i_1 
       (.I0(text[17]),
        .I1(cipher[49]),
        .I2(ready),
        .O(p_0_in[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair11" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[18]_i_1 
       (.I0(text[18]),
        .I1(cipher[50]),
        .I2(ready),
        .O(p_0_in[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair12" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[19]_i_1 
       (.I0(text[19]),
        .I1(cipher[51]),
        .I2(ready),
        .O(p_0_in[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair1" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[1]_i_1 
       (.I0(text[1]),
        .I1(cipher[33]),
        .I2(ready),
        .O(p_0_in[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[20]_i_1 
       (.I0(text[20]),
        .I1(cipher[52]),
        .I2(ready),
        .O(p_0_in[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[21]_i_1 
       (.I0(text[21]),
        .I1(cipher[53]),
        .I2(ready),
        .O(p_0_in[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[22]_i_1 
       (.I0(text[22]),
        .I1(cipher[54]),
        .I2(ready),
        .O(p_0_in[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[23]_i_1 
       (.I0(text[23]),
        .I1(cipher[55]),
        .I2(ready),
        .O(p_0_in[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair15" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[24]_i_1 
       (.I0(text[24]),
        .I1(cipher[56]),
        .I2(ready),
        .O(p_0_in[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair15" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[25]_i_1 
       (.I0(text[25]),
        .I1(cipher[57]),
        .I2(ready),
        .O(p_0_in[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair16" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[26]_i_1 
       (.I0(text[26]),
        .I1(cipher[58]),
        .I2(ready),
        .O(p_0_in[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair16" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[27]_i_1 
       (.I0(text[27]),
        .I1(cipher[59]),
        .I2(ready),
        .O(p_0_in[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair17" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[28]_i_1 
       (.I0(text[28]),
        .I1(cipher[60]),
        .I2(ready),
        .O(p_0_in[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair17" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[29]_i_1 
       (.I0(text[29]),
        .I1(cipher[61]),
        .I2(ready),
        .O(p_0_in[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[2]_i_1 
       (.I0(text[2]),
        .I1(cipher[34]),
        .I2(ready),
        .O(p_0_in[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair18" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[30]_i_1 
       (.I0(text[30]),
        .I1(cipher[62]),
        .I2(ready),
        .O(p_0_in[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair18" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[31]_i_1 
       (.I0(text[31]),
        .I1(cipher[63]),
        .I2(ready),
        .O(p_0_in[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[3]_i_1 
       (.I0(text[3]),
        .I1(cipher[35]),
        .I2(ready),
        .O(p_0_in[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[4]_i_1 
       (.I0(text[4]),
        .I1(cipher[36]),
        .I2(ready),
        .O(p_0_in[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[5]_i_1 
       (.I0(text[5]),
        .I1(cipher[37]),
        .I2(ready),
        .O(p_0_in[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[6]_i_1 
       (.I0(text[6]),
        .I1(cipher[38]),
        .I2(ready),
        .O(p_0_in[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[7]_i_1 
       (.I0(text[7]),
        .I1(cipher[39]),
        .I2(ready),
        .O(p_0_in[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[8]_i_1 
       (.I0(text[8]),
        .I1(cipher[40]),
        .I2(ready),
        .O(p_0_in[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v0[9]_i_1 
       (.I0(text[9]),
        .I1(cipher[41]),
        .I2(ready),
        .O(p_0_in[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[0] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[0]),
        .Q(cipher[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[10] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[10]),
        .Q(cipher[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[11] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[11]),
        .Q(cipher[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[12] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[12]),
        .Q(cipher[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[13] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[13]),
        .Q(cipher[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[14] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[14]),
        .Q(cipher[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[15] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[15]),
        .Q(cipher[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[16] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[16]),
        .Q(cipher[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[17] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[17]),
        .Q(cipher[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[18] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[18]),
        .Q(cipher[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[19] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[19]),
        .Q(cipher[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[1] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[1]),
        .Q(cipher[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[20] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[20]),
        .Q(cipher[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[21] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[21]),
        .Q(cipher[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[22] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[22]),
        .Q(cipher[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[23] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[23]),
        .Q(cipher[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[24] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[24]),
        .Q(cipher[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[25] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[25]),
        .Q(cipher[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[26] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[26]),
        .Q(cipher[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[27] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[27]),
        .Q(cipher[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[28] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[28]),
        .Q(cipher[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[29] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[29]),
        .Q(cipher[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[2] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[2]),
        .Q(cipher[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[30] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[30]),
        .Q(cipher[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[31] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[31]),
        .Q(cipher[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[3] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[3]),
        .Q(cipher[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[4] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[4]),
        .Q(cipher[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[5] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[5]),
        .Q(cipher[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[6] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[6]),
        .Q(cipher[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[7] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[7]),
        .Q(cipher[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[8] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[8]),
        .Q(cipher[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v0_reg[9] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(p_0_in[9]),
        .Q(cipher[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[11]_i_13 
       (.I0(cipher[43]),
        .I1(sum_reg[11]),
        .O(v1));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[11]_i_14 
       (.I0(cipher[42]),
        .I1(sum_reg[10]),
        .O(\v1[11]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[11]_i_15 
       (.I0(cipher[41]),
        .I1(sum_reg[9]),
        .O(\v1[11]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[11]_i_16 
       (.I0(cipher[40]),
        .I1(sum_reg[8]),
        .O(\v1[11]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[11]_i_17 
       (.I0(cipher[48]),
        .I1(sel),
        .I2(k1[11]),
        .I3(k3[11]),
        .O(\v1[11]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[11]_i_18 
       (.I0(cipher[47]),
        .I1(sel),
        .I2(k1[10]),
        .I3(k3[10]),
        .O(\v1[11]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[11]_i_19 
       (.I0(cipher[46]),
        .I1(sel),
        .I2(k1[9]),
        .I3(k3[9]),
        .O(\v1[11]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[11]_i_2 
       (.I0(plusOp0_out[11]),
        .I1(plusOp1_out[11]),
        .I2(plusOp[11]),
        .I3(ready),
        .O(\v1[11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[11]_i_20 
       (.I0(cipher[45]),
        .I1(sel),
        .I2(k1[8]),
        .I3(k3[8]),
        .O(\v1[11]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[11]_i_21 
       (.I0(cipher[38]),
        .I1(sel),
        .I2(k0[10]),
        .I3(k2[10]),
        .O(\v1[11]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[11]_i_22 
       (.I0(cipher[37]),
        .I1(sel),
        .I2(k0[9]),
        .I3(k2[9]),
        .O(\v1[11]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[11]_i_23 
       (.I0(cipher[36]),
        .I1(sel),
        .I2(k0[8]),
        .I3(k2[8]),
        .O(\v1[11]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[11]_i_24 
       (.I0(cipher[35]),
        .I1(sel),
        .I2(k0[7]),
        .I3(k2[7]),
        .O(\v1[11]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[11]_i_3 
       (.I0(plusOp0_out[10]),
        .I1(plusOp1_out[10]),
        .I2(plusOp[10]),
        .I3(ready),
        .O(\v1[11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[11]_i_4 
       (.I0(plusOp0_out[9]),
        .I1(plusOp1_out[9]),
        .I2(plusOp[9]),
        .I3(ready),
        .O(\v1[11]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[11]_i_5 
       (.I0(plusOp0_out[8]),
        .I1(plusOp1_out[8]),
        .I2(plusOp[8]),
        .I3(ready),
        .O(\v1[11]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[11]_i_6 
       (.I0(plusOp[11]),
        .I1(plusOp1_out[11]),
        .I2(plusOp0_out[11]),
        .I3(cipher[11]),
        .I4(ready),
        .I5(text[43]),
        .O(\v1[11]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[11]_i_7 
       (.I0(plusOp[10]),
        .I1(plusOp1_out[10]),
        .I2(plusOp0_out[10]),
        .I3(cipher[10]),
        .I4(ready),
        .I5(text[42]),
        .O(\v1[11]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[11]_i_8 
       (.I0(plusOp[9]),
        .I1(plusOp1_out[9]),
        .I2(plusOp0_out[9]),
        .I3(cipher[9]),
        .I4(ready),
        .I5(text[41]),
        .O(\v1[11]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[11]_i_9 
       (.I0(plusOp[8]),
        .I1(plusOp1_out[8]),
        .I2(plusOp0_out[8]),
        .I3(cipher[8]),
        .I4(ready),
        .I5(text[40]),
        .O(\v1[11]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[15]_i_13 
       (.I0(cipher[47]),
        .I1(sum_reg[15]),
        .O(\v1[15]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[15]_i_14 
       (.I0(cipher[46]),
        .I1(sum_reg[14]),
        .O(\v1[15]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[15]_i_15 
       (.I0(cipher[45]),
        .I1(sum_reg[13]),
        .O(\v1[15]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[15]_i_16 
       (.I0(cipher[44]),
        .I1(sum_reg[12]),
        .O(\v1[15]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[15]_i_17 
       (.I0(cipher[52]),
        .I1(sel),
        .I2(k1[15]),
        .I3(k3[15]),
        .O(\v1[15]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[15]_i_18 
       (.I0(cipher[51]),
        .I1(sel),
        .I2(k1[14]),
        .I3(k3[14]),
        .O(\v1[15]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[15]_i_19 
       (.I0(cipher[50]),
        .I1(sel),
        .I2(k1[13]),
        .I3(k3[13]),
        .O(\v1[15]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[15]_i_2 
       (.I0(plusOp0_out[15]),
        .I1(plusOp1_out[15]),
        .I2(plusOp[15]),
        .I3(ready),
        .O(\v1[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[15]_i_20 
       (.I0(cipher[49]),
        .I1(sel),
        .I2(k1[12]),
        .I3(k3[12]),
        .O(\v1[15]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[15]_i_21 
       (.I0(cipher[42]),
        .I1(sel),
        .I2(k0[14]),
        .I3(k2[14]),
        .O(\v1[15]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[15]_i_22 
       (.I0(cipher[41]),
        .I1(sel),
        .I2(k0[13]),
        .I3(k2[13]),
        .O(\v1[15]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[15]_i_23 
       (.I0(cipher[40]),
        .I1(sel),
        .I2(k0[12]),
        .I3(k2[12]),
        .O(\v1[15]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[15]_i_24 
       (.I0(cipher[39]),
        .I1(sel),
        .I2(k0[11]),
        .I3(k2[11]),
        .O(\v1[15]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[15]_i_3 
       (.I0(plusOp0_out[14]),
        .I1(plusOp1_out[14]),
        .I2(plusOp[14]),
        .I3(ready),
        .O(\v1[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[15]_i_4 
       (.I0(plusOp0_out[13]),
        .I1(plusOp1_out[13]),
        .I2(plusOp[13]),
        .I3(ready),
        .O(\v1[15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[15]_i_5 
       (.I0(plusOp0_out[12]),
        .I1(plusOp1_out[12]),
        .I2(plusOp[12]),
        .I3(ready),
        .O(\v1[15]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[15]_i_6 
       (.I0(plusOp[15]),
        .I1(plusOp1_out[15]),
        .I2(plusOp0_out[15]),
        .I3(cipher[15]),
        .I4(ready),
        .I5(text[47]),
        .O(\v1[15]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[15]_i_7 
       (.I0(plusOp[14]),
        .I1(plusOp1_out[14]),
        .I2(plusOp0_out[14]),
        .I3(cipher[14]),
        .I4(ready),
        .I5(text[46]),
        .O(\v1[15]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[15]_i_8 
       (.I0(plusOp[13]),
        .I1(plusOp1_out[13]),
        .I2(plusOp0_out[13]),
        .I3(cipher[13]),
        .I4(ready),
        .I5(text[45]),
        .O(\v1[15]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[15]_i_9 
       (.I0(plusOp[12]),
        .I1(plusOp1_out[12]),
        .I2(plusOp0_out[12]),
        .I3(cipher[12]),
        .I4(ready),
        .I5(text[44]),
        .O(\v1[15]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[19]_i_13 
       (.I0(cipher[51]),
        .I1(sum_reg[19]),
        .O(\v1[19]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[19]_i_14 
       (.I0(cipher[50]),
        .I1(sum_reg[18]),
        .O(\v1[19]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[19]_i_15 
       (.I0(cipher[49]),
        .I1(sum_reg[17]),
        .O(\v1[19]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[19]_i_16 
       (.I0(cipher[48]),
        .I1(sum_reg[16]),
        .O(\v1[19]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[19]_i_17 
       (.I0(cipher[56]),
        .I1(sel),
        .I2(k1[19]),
        .I3(k3[19]),
        .O(\v1[19]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[19]_i_18 
       (.I0(cipher[55]),
        .I1(sel),
        .I2(k1[18]),
        .I3(k3[18]),
        .O(\v1[19]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[19]_i_19 
       (.I0(cipher[54]),
        .I1(sel),
        .I2(k1[17]),
        .I3(k3[17]),
        .O(\v1[19]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[19]_i_2 
       (.I0(plusOp0_out[19]),
        .I1(plusOp1_out[19]),
        .I2(plusOp[19]),
        .I3(ready),
        .O(\v1[19]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[19]_i_20 
       (.I0(cipher[53]),
        .I1(sel),
        .I2(k1[16]),
        .I3(k3[16]),
        .O(\v1[19]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[19]_i_21 
       (.I0(cipher[46]),
        .I1(sel),
        .I2(k0[18]),
        .I3(k2[18]),
        .O(\v1[19]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[19]_i_22 
       (.I0(cipher[45]),
        .I1(sel),
        .I2(k0[17]),
        .I3(k2[17]),
        .O(\v1[19]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[19]_i_23 
       (.I0(cipher[44]),
        .I1(sel),
        .I2(k0[16]),
        .I3(k2[16]),
        .O(\v1[19]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[19]_i_24 
       (.I0(cipher[43]),
        .I1(sel),
        .I2(k0[15]),
        .I3(k2[15]),
        .O(\v1[19]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[19]_i_3 
       (.I0(plusOp0_out[18]),
        .I1(plusOp1_out[18]),
        .I2(plusOp[18]),
        .I3(ready),
        .O(\v1[19]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[19]_i_4 
       (.I0(plusOp0_out[17]),
        .I1(plusOp1_out[17]),
        .I2(plusOp[17]),
        .I3(ready),
        .O(\v1[19]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[19]_i_5 
       (.I0(plusOp0_out[16]),
        .I1(plusOp1_out[16]),
        .I2(plusOp[16]),
        .I3(ready),
        .O(\v1[19]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[19]_i_6 
       (.I0(plusOp[19]),
        .I1(plusOp1_out[19]),
        .I2(plusOp0_out[19]),
        .I3(cipher[19]),
        .I4(ready),
        .I5(text[51]),
        .O(\v1[19]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[19]_i_7 
       (.I0(plusOp[18]),
        .I1(plusOp1_out[18]),
        .I2(plusOp0_out[18]),
        .I3(cipher[18]),
        .I4(ready),
        .I5(text[50]),
        .O(\v1[19]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[19]_i_8 
       (.I0(plusOp[17]),
        .I1(plusOp1_out[17]),
        .I2(plusOp0_out[17]),
        .I3(cipher[17]),
        .I4(ready),
        .I5(text[49]),
        .O(\v1[19]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[19]_i_9 
       (.I0(plusOp[16]),
        .I1(plusOp1_out[16]),
        .I2(plusOp0_out[16]),
        .I3(cipher[16]),
        .I4(ready),
        .I5(text[48]),
        .O(\v1[19]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[23]_i_13 
       (.I0(cipher[55]),
        .I1(sum_reg[23]),
        .O(\v1[23]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[23]_i_14 
       (.I0(cipher[54]),
        .I1(sum_reg[22]),
        .O(\v1[23]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[23]_i_15 
       (.I0(cipher[53]),
        .I1(sum_reg[21]),
        .O(\v1[23]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[23]_i_16 
       (.I0(cipher[52]),
        .I1(sum_reg[20]),
        .O(\v1[23]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[23]_i_17 
       (.I0(cipher[60]),
        .I1(sel),
        .I2(k1[23]),
        .I3(k3[23]),
        .O(\v1[23]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[23]_i_18 
       (.I0(cipher[59]),
        .I1(sel),
        .I2(k1[22]),
        .I3(k3[22]),
        .O(\v1[23]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[23]_i_19 
       (.I0(cipher[58]),
        .I1(sel),
        .I2(k1[21]),
        .I3(k3[21]),
        .O(\v1[23]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[23]_i_2 
       (.I0(plusOp0_out[23]),
        .I1(plusOp1_out[23]),
        .I2(plusOp[23]),
        .I3(ready),
        .O(\v1[23]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[23]_i_20 
       (.I0(cipher[57]),
        .I1(sel),
        .I2(k1[20]),
        .I3(k3[20]),
        .O(\v1[23]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[23]_i_21 
       (.I0(cipher[50]),
        .I1(sel),
        .I2(k0[22]),
        .I3(k2[22]),
        .O(\v1[23]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[23]_i_22 
       (.I0(cipher[49]),
        .I1(sel),
        .I2(k0[21]),
        .I3(k2[21]),
        .O(\v1[23]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[23]_i_23 
       (.I0(cipher[48]),
        .I1(sel),
        .I2(k0[20]),
        .I3(k2[20]),
        .O(\v1[23]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[23]_i_24 
       (.I0(cipher[47]),
        .I1(sel),
        .I2(k0[19]),
        .I3(k2[19]),
        .O(\v1[23]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[23]_i_3 
       (.I0(plusOp0_out[22]),
        .I1(plusOp1_out[22]),
        .I2(plusOp[22]),
        .I3(ready),
        .O(\v1[23]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[23]_i_4 
       (.I0(plusOp0_out[21]),
        .I1(plusOp1_out[21]),
        .I2(plusOp[21]),
        .I3(ready),
        .O(\v1[23]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[23]_i_5 
       (.I0(plusOp0_out[20]),
        .I1(plusOp1_out[20]),
        .I2(plusOp[20]),
        .I3(ready),
        .O(\v1[23]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[23]_i_6 
       (.I0(plusOp[23]),
        .I1(plusOp1_out[23]),
        .I2(plusOp0_out[23]),
        .I3(cipher[23]),
        .I4(ready),
        .I5(text[55]),
        .O(\v1[23]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[23]_i_7 
       (.I0(plusOp[22]),
        .I1(plusOp1_out[22]),
        .I2(plusOp0_out[22]),
        .I3(cipher[22]),
        .I4(ready),
        .I5(text[54]),
        .O(\v1[23]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[23]_i_8 
       (.I0(plusOp[21]),
        .I1(plusOp1_out[21]),
        .I2(plusOp0_out[21]),
        .I3(cipher[21]),
        .I4(ready),
        .I5(text[53]),
        .O(\v1[23]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[23]_i_9 
       (.I0(plusOp[20]),
        .I1(plusOp1_out[20]),
        .I2(plusOp0_out[20]),
        .I3(cipher[20]),
        .I4(ready),
        .I5(text[52]),
        .O(\v1[23]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[27]_i_13 
       (.I0(cipher[59]),
        .I1(sum_reg[27]),
        .O(\v1[27]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[27]_i_14 
       (.I0(cipher[58]),
        .I1(sum_reg[26]),
        .O(\v1[27]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[27]_i_15 
       (.I0(cipher[57]),
        .I1(sum_reg[25]),
        .O(\v1[27]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[27]_i_16 
       (.I0(cipher[56]),
        .I1(sum_reg[24]),
        .O(\v1[27]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v1[27]_i_17 
       (.I0(k3[27]),
        .I1(k1[27]),
        .I2(sel),
        .O(feistelKey1[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[27]_i_18 
       (.I0(cipher[63]),
        .I1(sel),
        .I2(k1[26]),
        .I3(k3[26]),
        .O(\v1[27]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[27]_i_19 
       (.I0(cipher[62]),
        .I1(sel),
        .I2(k1[25]),
        .I3(k3[25]),
        .O(\v1[27]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[27]_i_2 
       (.I0(plusOp0_out[27]),
        .I1(plusOp1_out[27]),
        .I2(plusOp[27]),
        .I3(ready),
        .O(\v1[27]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[27]_i_20 
       (.I0(cipher[61]),
        .I1(sel),
        .I2(k1[24]),
        .I3(k3[24]),
        .O(\v1[27]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[27]_i_21 
       (.I0(cipher[54]),
        .I1(sel),
        .I2(k0[26]),
        .I3(k2[26]),
        .O(\v1[27]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[27]_i_22 
       (.I0(cipher[53]),
        .I1(sel),
        .I2(k0[25]),
        .I3(k2[25]),
        .O(\v1[27]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[27]_i_23 
       (.I0(cipher[52]),
        .I1(sel),
        .I2(k0[24]),
        .I3(k2[24]),
        .O(\v1[27]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[27]_i_24 
       (.I0(cipher[51]),
        .I1(sel),
        .I2(k0[23]),
        .I3(k2[23]),
        .O(\v1[27]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[27]_i_3 
       (.I0(plusOp0_out[26]),
        .I1(plusOp1_out[26]),
        .I2(plusOp[26]),
        .I3(ready),
        .O(\v1[27]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[27]_i_4 
       (.I0(plusOp0_out[25]),
        .I1(plusOp1_out[25]),
        .I2(plusOp[25]),
        .I3(ready),
        .O(\v1[27]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[27]_i_5 
       (.I0(plusOp0_out[24]),
        .I1(plusOp1_out[24]),
        .I2(plusOp[24]),
        .I3(ready),
        .O(\v1[27]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[27]_i_6 
       (.I0(plusOp[27]),
        .I1(plusOp1_out[27]),
        .I2(plusOp0_out[27]),
        .I3(cipher[27]),
        .I4(ready),
        .I5(text[59]),
        .O(\v1[27]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[27]_i_7 
       (.I0(plusOp[26]),
        .I1(plusOp1_out[26]),
        .I2(plusOp0_out[26]),
        .I3(cipher[26]),
        .I4(ready),
        .I5(text[58]),
        .O(\v1[27]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[27]_i_8 
       (.I0(plusOp[25]),
        .I1(plusOp1_out[25]),
        .I2(plusOp0_out[25]),
        .I3(cipher[25]),
        .I4(ready),
        .I5(text[57]),
        .O(\v1[27]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[27]_i_9 
       (.I0(plusOp[24]),
        .I1(plusOp1_out[24]),
        .I2(plusOp0_out[24]),
        .I3(cipher[24]),
        .I4(ready),
        .I5(text[56]),
        .O(\v1[27]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[31]_i_13 
       (.I0(cipher[58]),
        .I1(sel),
        .I2(k0[30]),
        .I3(k2[30]),
        .O(\v1[31]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[31]_i_14 
       (.I0(cipher[57]),
        .I1(sel),
        .I2(k0[29]),
        .I3(k2[29]),
        .O(\v1[31]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[31]_i_15 
       (.I0(cipher[56]),
        .I1(sel),
        .I2(k0[28]),
        .I3(k2[28]),
        .O(\v1[31]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[31]_i_16 
       (.I0(cipher[55]),
        .I1(sel),
        .I2(k0[27]),
        .I3(k2[27]),
        .O(\v1[31]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[31]_i_17 
       (.I0(cipher[63]),
        .I1(sum_reg[31]),
        .O(\v1[31]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[31]_i_18 
       (.I0(cipher[62]),
        .I1(sum_reg[30]),
        .O(\v1[31]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[31]_i_19 
       (.I0(cipher[61]),
        .I1(sum_reg[29]),
        .O(\v1[31]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[31]_i_2 
       (.I0(plusOp0_out[30]),
        .I1(plusOp1_out[30]),
        .I2(plusOp[30]),
        .I3(ready),
        .O(\v1[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[31]_i_20 
       (.I0(cipher[60]),
        .I1(sum_reg[28]),
        .O(\v1[31]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v1[31]_i_21 
       (.I0(k3[31]),
        .I1(k1[31]),
        .I2(sel),
        .O(feistelKey1[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v1[31]_i_22 
       (.I0(k3[30]),
        .I1(k1[30]),
        .I2(sel),
        .O(feistelKey1[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v1[31]_i_23 
       (.I0(k3[29]),
        .I1(k1[29]),
        .I2(sel),
        .O(feistelKey1[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v1[31]_i_24 
       (.I0(k3[28]),
        .I1(k1[28]),
        .I2(sel),
        .O(feistelKey1[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[31]_i_25 
       (.I0(cipher[59]),
        .I1(sel),
        .I2(k0[31]),
        .I3(k2[31]),
        .O(\v1[31]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[31]_i_3 
       (.I0(plusOp0_out[29]),
        .I1(plusOp1_out[29]),
        .I2(plusOp[29]),
        .I3(ready),
        .O(\v1[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[31]_i_4 
       (.I0(plusOp0_out[28]),
        .I1(plusOp1_out[28]),
        .I2(plusOp[28]),
        .I3(ready),
        .O(\v1[31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[31]_i_5 
       (.I0(plusOp[31]),
        .I1(plusOp1_out[31]),
        .I2(plusOp0_out[31]),
        .I3(cipher[31]),
        .I4(ready),
        .I5(text[63]),
        .O(\v1[31]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[31]_i_6 
       (.I0(plusOp[30]),
        .I1(plusOp1_out[30]),
        .I2(plusOp0_out[30]),
        .I3(cipher[30]),
        .I4(ready),
        .I5(text[62]),
        .O(\v1[31]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[31]_i_7 
       (.I0(plusOp[29]),
        .I1(plusOp1_out[29]),
        .I2(plusOp0_out[29]),
        .I3(cipher[29]),
        .I4(ready),
        .I5(text[61]),
        .O(\v1[31]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[31]_i_8 
       (.I0(plusOp[28]),
        .I1(plusOp1_out[28]),
        .I2(plusOp0_out[28]),
        .I3(cipher[28]),
        .I4(ready),
        .I5(text[60]),
        .O(\v1[31]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v1[3]_i_12 
       (.I0(k2[2]),
        .I1(k0[2]),
        .I2(sel),
        .O(feistelKey0__0[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v1[3]_i_13 
       (.I0(k2[1]),
        .I1(k0[1]),
        .I2(sel),
        .O(feistelKey0__0[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v1[3]_i_14 
       (.I0(k2[0]),
        .I1(k0[0]),
        .I2(sel),
        .O(feistelKey0__0[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[3]_i_15 
       (.I0(cipher[35]),
        .I1(sum_reg[3]),
        .O(\v1[3]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[3]_i_16 
       (.I0(cipher[34]),
        .I1(sum_reg[2]),
        .O(\v1[3]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[3]_i_17 
       (.I0(cipher[33]),
        .I1(sum_reg[1]),
        .O(\v1[3]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[3]_i_18 
       (.I0(cipher[32]),
        .I1(sum_reg[0]),
        .O(\v1[3]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[3]_i_19 
       (.I0(cipher[40]),
        .I1(sel),
        .I2(k1[3]),
        .I3(k3[3]),
        .O(\v1[3]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[3]_i_2 
       (.I0(plusOp0_out[3]),
        .I1(plusOp1_out[3]),
        .I2(plusOp[3]),
        .I3(ready),
        .O(\v1[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[3]_i_20 
       (.I0(cipher[39]),
        .I1(sel),
        .I2(k1[2]),
        .I3(k3[2]),
        .O(\v1[3]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[3]_i_21 
       (.I0(cipher[38]),
        .I1(sel),
        .I2(k1[1]),
        .I3(k3[1]),
        .O(\v1[3]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[3]_i_22 
       (.I0(cipher[37]),
        .I1(sel),
        .I2(k1[0]),
        .I3(k3[0]),
        .O(\v1[3]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000AC5353AC)) 
    \v1[3]_i_3 
       (.I0(k2[2]),
        .I1(k0[2]),
        .I2(sel),
        .I3(plusOp1_out[2]),
        .I4(plusOp[2]),
        .I5(ready),
        .O(\v1[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000AC5353AC)) 
    \v1[3]_i_4 
       (.I0(k2[1]),
        .I1(k0[1]),
        .I2(sel),
        .I3(plusOp1_out[1]),
        .I4(plusOp[1]),
        .I5(ready),
        .O(\v1[3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000AC5353AC)) 
    \v1[3]_i_5 
       (.I0(k2[0]),
        .I1(k0[0]),
        .I2(sel),
        .I3(plusOp1_out[0]),
        .I4(plusOp[0]),
        .I5(ready),
        .O(\v1[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[3]_i_6 
       (.I0(plusOp[3]),
        .I1(plusOp1_out[3]),
        .I2(plusOp0_out[3]),
        .I3(cipher[3]),
        .I4(ready),
        .I5(text[35]),
        .O(\v1[3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[3]_i_7 
       (.I0(plusOp[2]),
        .I1(plusOp1_out[2]),
        .I2(feistelKey0__0[2]),
        .I3(cipher[2]),
        .I4(ready),
        .I5(text[34]),
        .O(\v1[3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[3]_i_8 
       (.I0(plusOp[1]),
        .I1(plusOp1_out[1]),
        .I2(feistelKey0__0[1]),
        .I3(cipher[1]),
        .I4(ready),
        .I5(text[33]),
        .O(\v1[3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[3]_i_9 
       (.I0(plusOp[0]),
        .I1(plusOp1_out[0]),
        .I2(feistelKey0__0[0]),
        .I3(cipher[0]),
        .I4(ready),
        .I5(text[32]),
        .O(\v1[3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[7]_i_13 
       (.I0(cipher[39]),
        .I1(sum_reg[7]),
        .O(\v1[7]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[7]_i_14 
       (.I0(cipher[38]),
        .I1(sum_reg[6]),
        .O(\v1[7]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[7]_i_15 
       (.I0(cipher[37]),
        .I1(sum_reg[5]),
        .O(\v1[7]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \v1[7]_i_16 
       (.I0(cipher[36]),
        .I1(sum_reg[4]),
        .O(\v1[7]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[7]_i_17 
       (.I0(cipher[44]),
        .I1(sel),
        .I2(k1[7]),
        .I3(k3[7]),
        .O(\v1[7]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[7]_i_18 
       (.I0(cipher[43]),
        .I1(sel),
        .I2(k1[6]),
        .I3(k3[6]),
        .O(\v1[7]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[7]_i_19 
       (.I0(cipher[42]),
        .I1(sel),
        .I2(k1[5]),
        .I3(k3[5]),
        .O(\v1[7]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[7]_i_2 
       (.I0(plusOp0_out[7]),
        .I1(plusOp1_out[7]),
        .I2(plusOp[7]),
        .I3(ready),
        .O(\v1[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[7]_i_20 
       (.I0(cipher[41]),
        .I1(sel),
        .I2(k1[4]),
        .I3(k3[4]),
        .O(\v1[7]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[7]_i_21 
       (.I0(cipher[34]),
        .I1(sel),
        .I2(k0[6]),
        .I3(k2[6]),
        .O(\v1[7]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[7]_i_22 
       (.I0(cipher[33]),
        .I1(sel),
        .I2(k0[5]),
        .I3(k2[5]),
        .O(\v1[7]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    \v1[7]_i_23 
       (.I0(cipher[32]),
        .I1(sel),
        .I2(k0[4]),
        .I3(k2[4]),
        .O(\v1[7]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \v1[7]_i_24 
       (.I0(k2[3]),
        .I1(k0[3]),
        .I2(sel),
        .O(feistelKey0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[7]_i_3 
       (.I0(plusOp0_out[6]),
        .I1(plusOp1_out[6]),
        .I2(plusOp[6]),
        .I3(ready),
        .O(\v1[7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[7]_i_4 
       (.I0(plusOp0_out[5]),
        .I1(plusOp1_out[5]),
        .I2(plusOp[5]),
        .I3(ready),
        .O(\v1[7]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0096)) 
    \v1[7]_i_5 
       (.I0(plusOp0_out[4]),
        .I1(plusOp1_out[4]),
        .I2(plusOp[4]),
        .I3(ready),
        .O(\v1[7]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[7]_i_6 
       (.I0(plusOp[7]),
        .I1(plusOp1_out[7]),
        .I2(plusOp0_out[7]),
        .I3(cipher[7]),
        .I4(ready),
        .I5(text[39]),
        .O(\v1[7]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[7]_i_7 
       (.I0(plusOp[6]),
        .I1(plusOp1_out[6]),
        .I2(plusOp0_out[6]),
        .I3(cipher[6]),
        .I4(ready),
        .I5(text[38]),
        .O(\v1[7]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[7]_i_8 
       (.I0(plusOp[5]),
        .I1(plusOp1_out[5]),
        .I2(plusOp0_out[5]),
        .I3(cipher[5]),
        .I4(ready),
        .I5(text[37]),
        .O(\v1[7]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF699600006996)) 
    \v1[7]_i_9 
       (.I0(plusOp[4]),
        .I1(plusOp1_out[4]),
        .I2(plusOp0_out[4]),
        .I3(cipher[4]),
        .I4(ready),
        .I5(text[36]),
        .O(\v1[7]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[0] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[3]_i_1_n_7 ),
        .Q(cipher[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[10] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[11]_i_1_n_5 ),
        .Q(cipher[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[11] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[11]_i_1_n_4 ),
        .Q(cipher[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[11]_i_1 
       (.CI(\v1_reg[7]_i_1_n_0 ),
        .CO({\v1_reg[11]_i_1_n_0 ,\v1_reg[11]_i_1_n_1 ,\v1_reg[11]_i_1_n_2 ,\v1_reg[11]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\v1[11]_i_2_n_0 ,\v1[11]_i_3_n_0 ,\v1[11]_i_4_n_0 ,\v1[11]_i_5_n_0 }),
        .O({\v1_reg[11]_i_1_n_4 ,\v1_reg[11]_i_1_n_5 ,\v1_reg[11]_i_1_n_6 ,\v1_reg[11]_i_1_n_7 }),
        .S({\v1[11]_i_6_n_0 ,\v1[11]_i_7_n_0 ,\v1[11]_i_8_n_0 ,\v1[11]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[11]_i_10 
       (.CI(\v1_reg[7]_i_10_n_0 ),
        .CO(v1_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI(cipher[43:40]),
        .O(plusOp1_out[11:8]),
        .S({v1,\v1[11]_i_14_n_0 ,\v1[11]_i_15_n_0 ,\v1[11]_i_16_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[11]_i_11 
       (.CI(\v1_reg[7]_i_11_n_0 ),
        .CO({\v1_reg[11]_i_11_n_0 ,\v1_reg[11]_i_11_n_1 ,\v1_reg[11]_i_11_n_2 ,\v1_reg[11]_i_11_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(cipher[48:45]),
        .O(plusOp[11:8]),
        .S({\v1[11]_i_17_n_0 ,\v1[11]_i_18_n_0 ,\v1[11]_i_19_n_0 ,\v1[11]_i_20_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[11]_i_12 
       (.CI(\v1_reg[7]_i_12_n_0 ),
        .CO({\v1_reg[11]_i_12_n_0 ,\v1_reg[11]_i_12_n_1 ,\v1_reg[11]_i_12_n_2 ,\v1_reg[11]_i_12_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(cipher[38:35]),
        .O(plusOp0_out[10:7]),
        .S({\v1[11]_i_21_n_0 ,\v1[11]_i_22_n_0 ,\v1[11]_i_23_n_0 ,\v1[11]_i_24_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[12] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[15]_i_1_n_7 ),
        .Q(cipher[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[13] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[15]_i_1_n_6 ),
        .Q(cipher[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[14] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[15]_i_1_n_5 ),
        .Q(cipher[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[15] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[15]_i_1_n_4 ),
        .Q(cipher[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[15]_i_1 
       (.CI(\v1_reg[11]_i_1_n_0 ),
        .CO({\v1_reg[15]_i_1_n_0 ,\v1_reg[15]_i_1_n_1 ,\v1_reg[15]_i_1_n_2 ,\v1_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\v1[15]_i_2_n_0 ,\v1[15]_i_3_n_0 ,\v1[15]_i_4_n_0 ,\v1[15]_i_5_n_0 }),
        .O({\v1_reg[15]_i_1_n_4 ,\v1_reg[15]_i_1_n_5 ,\v1_reg[15]_i_1_n_6 ,\v1_reg[15]_i_1_n_7 }),
        .S({\v1[15]_i_6_n_0 ,\v1[15]_i_7_n_0 ,\v1[15]_i_8_n_0 ,\v1[15]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[15]_i_10 
       (.CI(v1_reg[3]),
        .CO({\v1_reg[15]_i_10_n_0 ,\v1_reg[15]_i_10_n_1 ,\v1_reg[15]_i_10_n_2 ,\v1_reg[15]_i_10_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(cipher[47:44]),
        .O(plusOp1_out[15:12]),
        .S({\v1[15]_i_13_n_0 ,\v1[15]_i_14_n_0 ,\v1[15]_i_15_n_0 ,\v1[15]_i_16_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[15]_i_11 
       (.CI(\v1_reg[11]_i_11_n_0 ),
        .CO({\v1_reg[15]_i_11_n_0 ,\v1_reg[15]_i_11_n_1 ,\v1_reg[15]_i_11_n_2 ,\v1_reg[15]_i_11_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(cipher[52:49]),
        .O(plusOp[15:12]),
        .S({\v1[15]_i_17_n_0 ,\v1[15]_i_18_n_0 ,\v1[15]_i_19_n_0 ,\v1[15]_i_20_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[15]_i_12 
       (.CI(\v1_reg[11]_i_12_n_0 ),
        .CO({\v1_reg[15]_i_12_n_0 ,\v1_reg[15]_i_12_n_1 ,\v1_reg[15]_i_12_n_2 ,\v1_reg[15]_i_12_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(cipher[42:39]),
        .O(plusOp0_out[14:11]),
        .S({\v1[15]_i_21_n_0 ,\v1[15]_i_22_n_0 ,\v1[15]_i_23_n_0 ,\v1[15]_i_24_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[16] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[19]_i_1_n_7 ),
        .Q(cipher[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[17] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[19]_i_1_n_6 ),
        .Q(cipher[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[18] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[19]_i_1_n_5 ),
        .Q(cipher[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[19] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[19]_i_1_n_4 ),
        .Q(cipher[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[19]_i_1 
       (.CI(\v1_reg[15]_i_1_n_0 ),
        .CO({\v1_reg[19]_i_1_n_0 ,\v1_reg[19]_i_1_n_1 ,\v1_reg[19]_i_1_n_2 ,\v1_reg[19]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\v1[19]_i_2_n_0 ,\v1[19]_i_3_n_0 ,\v1[19]_i_4_n_0 ,\v1[19]_i_5_n_0 }),
        .O({\v1_reg[19]_i_1_n_4 ,\v1_reg[19]_i_1_n_5 ,\v1_reg[19]_i_1_n_6 ,\v1_reg[19]_i_1_n_7 }),
        .S({\v1[19]_i_6_n_0 ,\v1[19]_i_7_n_0 ,\v1[19]_i_8_n_0 ,\v1[19]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[19]_i_10 
       (.CI(\v1_reg[15]_i_10_n_0 ),
        .CO({\v1_reg[19]_i_10_n_0 ,\v1_reg[19]_i_10_n_1 ,\v1_reg[19]_i_10_n_2 ,\v1_reg[19]_i_10_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(cipher[51:48]),
        .O(plusOp1_out[19:16]),
        .S({\v1[19]_i_13_n_0 ,\v1[19]_i_14_n_0 ,\v1[19]_i_15_n_0 ,\v1[19]_i_16_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[19]_i_11 
       (.CI(\v1_reg[15]_i_11_n_0 ),
        .CO({\v1_reg[19]_i_11_n_0 ,\v1_reg[19]_i_11_n_1 ,\v1_reg[19]_i_11_n_2 ,\v1_reg[19]_i_11_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(cipher[56:53]),
        .O(plusOp[19:16]),
        .S({\v1[19]_i_17_n_0 ,\v1[19]_i_18_n_0 ,\v1[19]_i_19_n_0 ,\v1[19]_i_20_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[19]_i_12 
       (.CI(\v1_reg[15]_i_12_n_0 ),
        .CO({\v1_reg[19]_i_12_n_0 ,\v1_reg[19]_i_12_n_1 ,\v1_reg[19]_i_12_n_2 ,\v1_reg[19]_i_12_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(cipher[46:43]),
        .O(plusOp0_out[18:15]),
        .S({\v1[19]_i_21_n_0 ,\v1[19]_i_22_n_0 ,\v1[19]_i_23_n_0 ,\v1[19]_i_24_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[1] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[3]_i_1_n_6 ),
        .Q(cipher[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[20] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[23]_i_1_n_7 ),
        .Q(cipher[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[21] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[23]_i_1_n_6 ),
        .Q(cipher[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[22] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[23]_i_1_n_5 ),
        .Q(cipher[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[23] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[23]_i_1_n_4 ),
        .Q(cipher[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[23]_i_1 
       (.CI(\v1_reg[19]_i_1_n_0 ),
        .CO({\v1_reg[23]_i_1_n_0 ,\v1_reg[23]_i_1_n_1 ,\v1_reg[23]_i_1_n_2 ,\v1_reg[23]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\v1[23]_i_2_n_0 ,\v1[23]_i_3_n_0 ,\v1[23]_i_4_n_0 ,\v1[23]_i_5_n_0 }),
        .O({\v1_reg[23]_i_1_n_4 ,\v1_reg[23]_i_1_n_5 ,\v1_reg[23]_i_1_n_6 ,\v1_reg[23]_i_1_n_7 }),
        .S({\v1[23]_i_6_n_0 ,\v1[23]_i_7_n_0 ,\v1[23]_i_8_n_0 ,\v1[23]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[23]_i_10 
       (.CI(\v1_reg[19]_i_10_n_0 ),
        .CO({\v1_reg[23]_i_10_n_0 ,\v1_reg[23]_i_10_n_1 ,\v1_reg[23]_i_10_n_2 ,\v1_reg[23]_i_10_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(cipher[55:52]),
        .O(plusOp1_out[23:20]),
        .S({\v1[23]_i_13_n_0 ,\v1[23]_i_14_n_0 ,\v1[23]_i_15_n_0 ,\v1[23]_i_16_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[23]_i_11 
       (.CI(\v1_reg[19]_i_11_n_0 ),
        .CO({\v1_reg[23]_i_11_n_0 ,\v1_reg[23]_i_11_n_1 ,\v1_reg[23]_i_11_n_2 ,\v1_reg[23]_i_11_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(cipher[60:57]),
        .O(plusOp[23:20]),
        .S({\v1[23]_i_17_n_0 ,\v1[23]_i_18_n_0 ,\v1[23]_i_19_n_0 ,\v1[23]_i_20_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[23]_i_12 
       (.CI(\v1_reg[19]_i_12_n_0 ),
        .CO({\v1_reg[23]_i_12_n_0 ,\v1_reg[23]_i_12_n_1 ,\v1_reg[23]_i_12_n_2 ,\v1_reg[23]_i_12_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(cipher[50:47]),
        .O(plusOp0_out[22:19]),
        .S({\v1[23]_i_21_n_0 ,\v1[23]_i_22_n_0 ,\v1[23]_i_23_n_0 ,\v1[23]_i_24_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[24] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[27]_i_1_n_7 ),
        .Q(cipher[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[25] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[27]_i_1_n_6 ),
        .Q(cipher[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[26] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[27]_i_1_n_5 ),
        .Q(cipher[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[27] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[27]_i_1_n_4 ),
        .Q(cipher[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[27]_i_1 
       (.CI(\v1_reg[23]_i_1_n_0 ),
        .CO({\v1_reg[27]_i_1_n_0 ,\v1_reg[27]_i_1_n_1 ,\v1_reg[27]_i_1_n_2 ,\v1_reg[27]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\v1[27]_i_2_n_0 ,\v1[27]_i_3_n_0 ,\v1[27]_i_4_n_0 ,\v1[27]_i_5_n_0 }),
        .O({\v1_reg[27]_i_1_n_4 ,\v1_reg[27]_i_1_n_5 ,\v1_reg[27]_i_1_n_6 ,\v1_reg[27]_i_1_n_7 }),
        .S({\v1[27]_i_6_n_0 ,\v1[27]_i_7_n_0 ,\v1[27]_i_8_n_0 ,\v1[27]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[27]_i_10 
       (.CI(\v1_reg[23]_i_10_n_0 ),
        .CO({\v1_reg[27]_i_10_n_0 ,\v1_reg[27]_i_10_n_1 ,\v1_reg[27]_i_10_n_2 ,\v1_reg[27]_i_10_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(cipher[59:56]),
        .O(plusOp1_out[27:24]),
        .S({\v1[27]_i_13_n_0 ,\v1[27]_i_14_n_0 ,\v1[27]_i_15_n_0 ,\v1[27]_i_16_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[27]_i_11 
       (.CI(\v1_reg[23]_i_11_n_0 ),
        .CO({\v1_reg[27]_i_11_n_0 ,\v1_reg[27]_i_11_n_1 ,\v1_reg[27]_i_11_n_2 ,\v1_reg[27]_i_11_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,cipher[63:61]}),
        .O(plusOp[27:24]),
        .S({feistelKey1[27],\v1[27]_i_18_n_0 ,\v1[27]_i_19_n_0 ,\v1[27]_i_20_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[27]_i_12 
       (.CI(\v1_reg[23]_i_12_n_0 ),
        .CO({\v1_reg[27]_i_12_n_0 ,\v1_reg[27]_i_12_n_1 ,\v1_reg[27]_i_12_n_2 ,\v1_reg[27]_i_12_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(cipher[54:51]),
        .O(plusOp0_out[26:23]),
        .S({\v1[27]_i_21_n_0 ,\v1[27]_i_22_n_0 ,\v1[27]_i_23_n_0 ,\v1[27]_i_24_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[28] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[31]_i_1_n_7 ),
        .Q(cipher[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[29] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[31]_i_1_n_6 ),
        .Q(cipher[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[2] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[3]_i_1_n_5 ),
        .Q(cipher[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[30] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[31]_i_1_n_5 ),
        .Q(cipher[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[31] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[31]_i_1_n_4 ),
        .Q(cipher[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[31]_i_1 
       (.CI(\v1_reg[27]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\v1[31]_i_2_n_0 ,\v1[31]_i_3_n_0 ,\v1[31]_i_4_n_0 }),
        .O({\v1_reg[31]_i_1_n_4 ,\v1_reg[31]_i_1_n_5 ,\v1_reg[31]_i_1_n_6 ,\v1_reg[31]_i_1_n_7 }),
        .S({\v1[31]_i_5_n_0 ,\v1[31]_i_6_n_0 ,\v1[31]_i_7_n_0 ,\v1[31]_i_8_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[31]_i_10 
       (.CI(\v1_reg[27]_i_10_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,cipher[62:60]}),
        .O(plusOp1_out[31:28]),
        .S({\v1[31]_i_17_n_0 ,\v1[31]_i_18_n_0 ,\v1[31]_i_19_n_0 ,\v1[31]_i_20_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[31]_i_11 
       (.CI(\v1_reg[27]_i_11_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(plusOp[31:28]),
        .S(feistelKey1[31:28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[31]_i_12 
       (.CI(\v1_reg[31]_i_9_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\v1_reg[31]_i_12_n_4 ,\v1_reg[31]_i_12_n_5 ,\v1_reg[31]_i_12_n_6 ,plusOp0_out[31]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\v1[31]_i_25_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[31]_i_9 
       (.CI(\v1_reg[27]_i_12_n_0 ),
        .CO({\v1_reg[31]_i_9_n_0 ,\v1_reg[31]_i_9_n_1 ,\v1_reg[31]_i_9_n_2 ,\v1_reg[31]_i_9_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(cipher[58:55]),
        .O(plusOp0_out[30:27]),
        .S({\v1[31]_i_13_n_0 ,\v1[31]_i_14_n_0 ,\v1[31]_i_15_n_0 ,\v1[31]_i_16_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[3] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[3]_i_1_n_4 ),
        .Q(cipher[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[3]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO({\v1_reg[3]_i_1_n_0 ,\v1_reg[3]_i_1_n_1 ,\v1_reg[3]_i_1_n_2 ,\v1_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\v1[3]_i_2_n_0 ,\v1[3]_i_3_n_0 ,\v1[3]_i_4_n_0 ,\v1[3]_i_5_n_0 }),
        .O({\v1_reg[3]_i_1_n_4 ,\v1_reg[3]_i_1_n_5 ,\v1_reg[3]_i_1_n_6 ,\v1_reg[3]_i_1_n_7 }),
        .S({\v1[3]_i_6_n_0 ,\v1[3]_i_7_n_0 ,\v1[3]_i_8_n_0 ,\v1[3]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[3]_i_10 
       (.CI(\<const0>__0__0 ),
        .CO({\v1_reg[3]_i_10_n_0 ,\v1_reg[3]_i_10_n_1 ,\v1_reg[3]_i_10_n_2 ,\v1_reg[3]_i_10_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(cipher[35:32]),
        .O(plusOp1_out[3:0]),
        .S({\v1[3]_i_15_n_0 ,\v1[3]_i_16_n_0 ,\v1[3]_i_17_n_0 ,\v1[3]_i_18_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[3]_i_11 
       (.CI(\<const0>__0__0 ),
        .CO({\v1_reg[3]_i_11_n_0 ,\v1_reg[3]_i_11_n_1 ,\v1_reg[3]_i_11_n_2 ,\v1_reg[3]_i_11_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(cipher[40:37]),
        .O(plusOp[3:0]),
        .S({\v1[3]_i_19_n_0 ,\v1[3]_i_20_n_0 ,\v1[3]_i_21_n_0 ,\v1[3]_i_22_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[4] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[7]_i_1_n_7 ),
        .Q(cipher[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[5] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[7]_i_1_n_6 ),
        .Q(cipher[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[6] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[7]_i_1_n_5 ),
        .Q(cipher[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[7] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[7]_i_1_n_4 ),
        .Q(cipher[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[7]_i_1 
       (.CI(\v1_reg[3]_i_1_n_0 ),
        .CO({\v1_reg[7]_i_1_n_0 ,\v1_reg[7]_i_1_n_1 ,\v1_reg[7]_i_1_n_2 ,\v1_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\v1[7]_i_2_n_0 ,\v1[7]_i_3_n_0 ,\v1[7]_i_4_n_0 ,\v1[7]_i_5_n_0 }),
        .O({\v1_reg[7]_i_1_n_4 ,\v1_reg[7]_i_1_n_5 ,\v1_reg[7]_i_1_n_6 ,\v1_reg[7]_i_1_n_7 }),
        .S({\v1[7]_i_6_n_0 ,\v1[7]_i_7_n_0 ,\v1[7]_i_8_n_0 ,\v1[7]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[7]_i_10 
       (.CI(\v1_reg[3]_i_10_n_0 ),
        .CO({\v1_reg[7]_i_10_n_0 ,\v1_reg[7]_i_10_n_1 ,\v1_reg[7]_i_10_n_2 ,\v1_reg[7]_i_10_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(cipher[39:36]),
        .O(plusOp1_out[7:4]),
        .S({\v1[7]_i_13_n_0 ,\v1[7]_i_14_n_0 ,\v1[7]_i_15_n_0 ,\v1[7]_i_16_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[7]_i_11 
       (.CI(\v1_reg[3]_i_11_n_0 ),
        .CO({\v1_reg[7]_i_11_n_0 ,\v1_reg[7]_i_11_n_1 ,\v1_reg[7]_i_11_n_2 ,\v1_reg[7]_i_11_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(cipher[44:41]),
        .O(plusOp[7:4]),
        .S({\v1[7]_i_17_n_0 ,\v1[7]_i_18_n_0 ,\v1[7]_i_19_n_0 ,\v1[7]_i_20_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \v1_reg[7]_i_12 
       (.CI(\<const0>__0__0 ),
        .CO({\v1_reg[7]_i_12_n_0 ,\v1_reg[7]_i_12_n_1 ,\v1_reg[7]_i_12_n_2 ,\v1_reg[7]_i_12_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({cipher[34:32],\<const0>__0__0 }),
        .O(plusOp0_out[6:3]),
        .S({\v1[7]_i_21_n_0 ,\v1[7]_i_22_n_0 ,\v1[7]_i_23_n_0 ,feistelKey0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[8] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[11]_i_1_n_7 ),
        .Q(cipher[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \v1_reg[9] 
       (.C(clock),
        .CE(\<const1>__0__0 ),
        .D(\v1_reg[11]_i_1_n_6 ),
        .Q(cipher[41]),
        .R(\<const0>__0__0 ));
endmodule
