module aes128
   (clk,
    state,
    key,
    backdoor,
    out);
  output backdoor;
  input clk;
  input [127:0]state;
  input [127:0]key;
  output [127:0]out;

  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const0>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const1>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_1/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_1/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_1/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_1/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_1/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_1/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_1/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_1/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_1/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_1/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_1/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_1/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_1/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_1/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_1/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_1/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_3/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_3/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_3/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_3/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_3/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_3/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_3/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_3/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_3/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_3/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_3/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_3/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_3/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_3/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_3/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/S4_0/S_3/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a1/k0a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a1/k1a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a1/k2a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a1/k3a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a1/k4a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a1/v0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a1/v1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a1/v2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a1/v3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_1/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_1/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_1/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_1/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_1/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_1/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_1/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_1/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_1/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_1/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_1/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_1/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_1/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_1/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_1/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_1/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_3/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_3/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_3/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_3/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_3/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_3/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_3/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_3/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_3/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_3/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_3/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_3/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_3/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_3/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_3/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a10/S4_0/S_3/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a10/k0a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a10/k1a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a10/k2a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a10/k3a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a10/k4a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [29:25]\a10/v0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a10/v1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a10/v2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a10/v3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_1/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_1/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_1/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_1/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_1/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_1/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_1/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_1/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_1/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_1/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_1/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_1/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_1/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_1/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_1/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_1/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_3/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_3/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_3/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_3/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_3/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_3/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_3/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_3/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_3/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_3/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_3/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_3/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_3/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_3/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_3/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/S4_0/S_3/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a2/k0a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a2/k1a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a2/k2a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a2/k3a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a2/k4a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a2/v0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a2/v1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a2/v2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a2/v3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_1/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_1/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_1/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_1/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_1/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_1/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_1/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_1/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_1/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_1/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_1/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_1/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_1/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_1/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_1/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_1/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_3/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_3/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_3/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_3/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_3/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_3/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_3/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_3/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_3/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_3/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_3/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_3/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_3/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_3/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_3/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/S4_0/S_3/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a3/k0a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a3/k1a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a3/k2a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a3/k3a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a3/k4a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a3/v0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a3/v1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a3/v2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a3/v3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_1/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_1/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_1/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_1/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_1/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_1/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_1/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_1/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_1/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_1/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_1/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_1/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_1/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_1/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_1/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_1/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_3/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_3/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_3/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_3/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_3/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_3/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_3/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_3/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_3/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_3/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_3/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_3/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_3/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_3/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_3/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/S4_0/S_3/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a4/k0a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a4/k1a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a4/k2a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a4/k3a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a4/k4a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a4/v0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a4/v1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a4/v2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a4/v3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_1/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_1/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_1/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_1/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_1/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_1/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_1/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_1/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_1/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_1/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_1/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_1/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_1/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_1/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_1/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_1/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_3/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_3/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_3/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_3/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_3/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_3/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_3/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_3/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_3/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_3/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_3/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_3/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_3/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_3/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_3/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/S4_0/S_3/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a5/k0a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a5/k1a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a5/k2a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a5/k3a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a5/k4a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a5/v0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a5/v1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a5/v2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a5/v3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_1/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_1/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_1/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_1/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_1/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_1/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_1/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_1/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_1/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_1/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_1/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_1/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_1/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_1/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_1/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_1/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_3/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_3/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_3/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_3/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_3/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_3/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_3/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_3/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_3/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_3/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_3/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_3/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_3/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_3/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_3/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/S4_0/S_3/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a6/k0a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a6/k1a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a6/k2a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a6/k3a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a6/k4a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a6/v0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a6/v1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a6/v2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a6/v3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_1/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_1/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_1/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_1/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_1/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_1/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_1/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_1/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_1/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_1/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_1/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_1/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_1/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_1/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_1/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_1/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_3/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_3/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_3/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_3/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_3/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_3/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_3/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_3/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_3/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_3/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_3/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_3/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_3/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_3/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_3/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/S4_0/S_3/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a7/k0a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a7/k1a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a7/k2a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a7/k3a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a7/k4a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a7/v0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a7/v1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a7/v2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a7/v3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_1/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_1/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_1/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_1/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_1/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_1/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_1/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_1/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_1/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_1/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_1/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_1/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_1/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_1/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_1/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_1/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_3/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_3/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_3/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_3/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_3/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_3/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_3/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_3/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_3/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_3/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_3/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_3/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_3/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_3/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_3/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/S4_0/S_3/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a8/k0a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a8/k1a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a8/k2a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a8/k3a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a8/k4a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a8/v0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [30:0]\a8/v1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a8/v2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a8/v3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_1/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_1/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_1/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_1/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_1/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_1/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_1/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_1/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_1/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_1/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_1/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_1/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_1/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_1/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_1/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_1/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_3/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_3/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_3/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_3/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_3/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_3/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_3/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_3/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_3/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_3/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_3/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_3/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_3/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_3/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_3/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9/S4_0/S_3/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a9/k0a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a9/k1a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a9/k2a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a9/k3a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a9/k4a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [28:24]\a9/v0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a9/v1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a9/v2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\a9/v3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire clk;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]k0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]k0b;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]k1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire k1a;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \k1a[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \k1a[25]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \k1a[25]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \k1a[25]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \k1a[26]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \k1a[26]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \k1a[27]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \k1a[27]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \k1a[28]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \k1a[28]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \k1a[28]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \k1a[29]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \k1a[29]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \k1a[30]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \k1a[31]_i_1__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]k1b;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]k2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]k2b;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]k3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]k3b;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]k4;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]k4b;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]k5;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]k5b;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]k6;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]k6b;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]k7;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]k7b;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]k8;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]k8b;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]k9;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]key;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]\r1/p_0_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t0/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t0/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t0/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t0/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t0/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t0/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t0/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t0/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t0/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t1/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t1/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t1/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t1/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t1/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t1/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t1/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t1/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t1/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t2/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t2/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t2/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t2/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t2/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t2/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t2/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t2/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t2/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t3/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t3/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t3/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t3/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t3/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t3/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r1/t3/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t3/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r1/t3/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]\r2/p_0_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t0/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t0/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t0/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t0/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t0/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t0/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t0/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t0/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t0/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t1/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t1/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t1/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t1/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t1/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t1/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t1/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t1/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t1/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t2/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t2/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t2/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t2/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t2/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t2/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t2/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t2/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t2/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t3/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t3/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t3/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t3/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t3/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t3/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r2/t3/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t3/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r2/t3/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]\r3/p_0_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t0/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t0/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t0/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t0/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t0/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t0/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t0/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t0/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t0/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t1/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t1/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t1/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t1/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t1/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t1/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t1/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t1/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t1/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t2/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t2/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t2/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t2/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t2/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t2/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t2/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t2/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t2/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t3/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t3/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t3/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t3/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t3/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t3/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r3/t3/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t3/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r3/t3/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]\r4/p_0_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t0/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t0/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t0/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t0/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t0/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t0/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t0/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t0/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t0/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t1/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t1/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t1/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t1/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t1/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t1/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t1/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t1/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t1/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t2/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t2/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t2/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t2/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t2/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t2/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t2/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t2/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t2/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t3/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t3/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t3/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t3/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t3/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t3/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r4/t3/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t3/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r4/t3/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]\r5/p_0_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t0/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t0/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t0/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t0/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t0/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t0/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t0/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t0/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t0/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t1/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t1/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t1/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t1/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t1/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t1/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t1/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t1/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t1/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t2/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t2/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t2/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t2/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t2/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t2/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t2/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t2/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t2/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t3/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t3/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t3/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t3/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t3/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t3/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r5/t3/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t3/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r5/t3/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]\r6/p_0_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t0/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t0/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t0/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t0/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t0/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t0/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t0/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t0/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t0/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t1/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t1/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t1/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t1/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t1/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t1/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t1/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t1/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t1/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t2/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t2/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t2/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t2/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t2/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t2/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t2/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t2/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t2/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t3/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t3/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t3/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t3/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t3/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t3/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r6/t3/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t3/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r6/t3/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]\r7/p_0_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t0/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t0/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t0/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t0/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t0/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t0/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t0/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t0/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t0/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t1/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t1/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t1/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t1/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t1/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t1/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t1/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t1/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t1/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t2/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t2/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t2/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t2/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t2/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t2/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t2/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t2/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t2/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t3/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t3/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t3/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t3/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t3/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t3/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r7/t3/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t3/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r7/t3/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]\r8/p_0_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t0/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t0/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t0/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t0/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t0/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t0/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t0/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t0/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t0/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t1/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t1/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t1/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t1/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t1/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t1/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t1/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t1/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t1/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t2/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t2/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t2/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t2/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t2/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t2/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t2/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t2/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t2/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t3/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t3/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t3/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t3/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t3/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t3/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r8/t3/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t3/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r8/t3/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]\r9/p_0_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t0/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t0/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t0/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t0/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t0/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t0/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t0/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t0/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t0/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t1/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t1/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t1/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t1/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t1/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t1/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t1/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t1/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t1/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t2/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t2/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t2/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t2/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t2/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t2/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t2/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t2/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t2/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t3/t0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t3/t0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t0/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t3/t1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t3/t1/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t3/t2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t3/t2/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s0/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s0/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s0/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s0/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s0/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s0/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s0/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s0/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s0/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s0/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s0/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s0/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s0/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s0/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s0/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s0/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s4/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s4/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s4/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s4/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s4/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s4/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s4/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s4/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s4/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s4/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s4/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s4/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s4/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s4/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s4/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r9/t3/t2/s4/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t3/t3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\r9/t3/t3/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_1/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_1/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_1/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_1/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_1/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_1/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_1/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_1/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_1/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_1/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_1/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_1/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_1/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_1/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_1/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_1/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_3/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_3/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_3/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_3/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_3/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_3/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_3/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_3/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_3/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_3/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_3/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_3/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_3/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_3/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_3/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_1/S_3/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_1/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_1/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_1/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_1/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_1/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_1/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_1/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_1/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_1/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_1/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_1/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_1/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_1/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_1/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_1/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_1/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_3/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_3/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_3/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_3/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_3/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_3/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_3/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_3/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_3/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_3/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_3/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_3/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_3/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_3/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_3/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_2/S_3/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_1/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_1/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_1/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_1/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_1/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_1/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_1/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_1/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_1/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_1/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_1/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_1/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_1/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_1/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_1/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_1/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_3/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_3/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_3/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_3/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_3/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_3/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_3/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_3/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_3/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_3/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_3/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_3/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_3/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_3/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_3/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_3/S_3/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_1/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_1/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_1/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_1/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_1/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_1/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_1/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_1/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_1/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_1/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_1/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_1/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_1/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_1/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_1/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_1/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_3/out_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_3/out_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_3/out_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_3/out_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_3/out_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_3/out_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_3/out_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_3/out_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_3/out_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_3/out_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_3/out_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_3/out_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_3/out_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_3/out_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_3/out_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rf/S4_4/S_3/out_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\rf/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\rf/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\rf/p_2_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\rf/p_3_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]\rf/p_4_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]s0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[100]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[101]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[102]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[103]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[104]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[105]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[106]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[107]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[108]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[109]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[110]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[111]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[112]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[113]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[114]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[115]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[116]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[117]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[118]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[119]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[120]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[121]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[122]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[123]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[124]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[125]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[126]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[127]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[18]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[22]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[26]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[30]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[32]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[33]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[34]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[35]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[36]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[37]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[38]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[39]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[40]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[41]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[42]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[43]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[44]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[45]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[46]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[47]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[48]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[49]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[50]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[51]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[52]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[53]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[54]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[55]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[56]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[57]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[58]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[59]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[60]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[61]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[62]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[63]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[64]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[65]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[66]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[67]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[68]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[69]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[70]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[71]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[72]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[73]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[74]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[75]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[76]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[77]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[78]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[79]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[80]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[81]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[82]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[83]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[84]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[85]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[86]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[87]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[88]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[89]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[90]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[91]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[92]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[93]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[94]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[95]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[96]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[97]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[98]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[99]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \s0[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]s1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]s2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]s3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]s4;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]s5;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]s6;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]s7;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]s8;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]s9;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]state;

  assign backdoor =  \rf/S4_4/S_3/out_reg_n_7  ;

  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND
       (.G(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC
       (.P(\<const1>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_0/S_1/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \a1/S4_0/S_1/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,k0[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,k0[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\a1/S4_0/S_1/out_reg_n_0 ,\a1/S4_0/S_1/out_reg_n_1 ,\a1/S4_0/S_1/out_reg_n_2 ,\a1/S4_0/S_1/out_reg_n_3 ,\a1/S4_0/S_1/out_reg_n_4 ,\a1/S4_0/S_1/out_reg_n_5 ,\a1/S4_0/S_1/out_reg_n_6 ,\a1/S4_0/S_1/out_reg_n_7 ,\a1/k4a [23:16]}),
        .DOBDO({\a1/S4_0/S_1/out_reg_n_16 ,\a1/S4_0/S_1/out_reg_n_17 ,\a1/S4_0/S_1/out_reg_n_18 ,\a1/S4_0/S_1/out_reg_n_19 ,\a1/S4_0/S_1/out_reg_n_20 ,\a1/S4_0/S_1/out_reg_n_21 ,\a1/S4_0/S_1/out_reg_n_22 ,\a1/S4_0/S_1/out_reg_n_23 ,\a1/k4a [31:24]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_0/S_3/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \a1/S4_0/S_3/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,k0[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,k0[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\a1/S4_0/S_3/out_reg_n_0 ,\a1/S4_0/S_3/out_reg_n_1 ,\a1/S4_0/S_3/out_reg_n_2 ,\a1/S4_0/S_3/out_reg_n_3 ,\a1/S4_0/S_3/out_reg_n_4 ,\a1/S4_0/S_3/out_reg_n_5 ,\a1/S4_0/S_3/out_reg_n_6 ,\a1/S4_0/S_3/out_reg_n_7 ,\a1/k4a [7:0]}),
        .DOBDO({\a1/S4_0/S_3/out_reg_n_16 ,\a1/S4_0/S_3/out_reg_n_17 ,\a1/S4_0/S_3/out_reg_n_18 ,\a1/S4_0/S_3/out_reg_n_19 ,\a1/S4_0/S_3/out_reg_n_20 ,\a1/S4_0/S_3/out_reg_n_21 ,\a1/S4_0/S_3/out_reg_n_22 ,\a1/S4_0/S_3/out_reg_n_23 ,\a1/k4a [15:8]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[96]),
        .Q(\a1/k0a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[106]),
        .Q(\a1/k0a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[107]),
        .Q(\a1/k0a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[108]),
        .Q(\a1/k0a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[109]),
        .Q(\a1/k0a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[110]),
        .Q(\a1/k0a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[111]),
        .Q(\a1/k0a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[112]),
        .Q(\a1/k0a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[113]),
        .Q(\a1/k0a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[114]),
        .Q(\a1/k0a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[115]),
        .Q(\a1/k0a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[97]),
        .Q(\a1/k0a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[116]),
        .Q(\a1/k0a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[117]),
        .Q(\a1/k0a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[118]),
        .Q(\a1/k0a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[119]),
        .Q(\a1/k0a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v0 ),
        .Q(\a1/k0a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[121]),
        .Q(\a1/k0a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[122]),
        .Q(\a1/k0a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[123]),
        .Q(\a1/k0a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[124]),
        .Q(\a1/k0a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[125]),
        .Q(\a1/k0a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[98]),
        .Q(\a1/k0a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[126]),
        .Q(\a1/k0a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[127]),
        .Q(\a1/k0a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[99]),
        .Q(\a1/k0a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[100]),
        .Q(\a1/k0a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[101]),
        .Q(\a1/k0a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[102]),
        .Q(\a1/k0a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[103]),
        .Q(\a1/k0a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[104]),
        .Q(\a1/k0a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k0a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0[105]),
        .Q(\a1/k0a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [0]),
        .Q(\a1/k1a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [10]),
        .Q(\a1/k1a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [11]),
        .Q(\a1/k1a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [12]),
        .Q(\a1/k1a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [13]),
        .Q(\a1/k1a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [14]),
        .Q(\a1/k1a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [15]),
        .Q(\a1/k1a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [16]),
        .Q(\a1/k1a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [17]),
        .Q(\a1/k1a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [18]),
        .Q(\a1/k1a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [19]),
        .Q(\a1/k1a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [1]),
        .Q(\a1/k1a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [20]),
        .Q(\a1/k1a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [21]),
        .Q(\a1/k1a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [22]),
        .Q(\a1/k1a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [23]),
        .Q(\a1/k1a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\k1a[24]_i_1_n_0 ),
        .Q(\a1/k1a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [25]),
        .Q(\a1/k1a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [26]),
        .Q(\a1/k1a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [27]),
        .Q(\a1/k1a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [28]),
        .Q(\a1/k1a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [29]),
        .Q(\a1/k1a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [2]),
        .Q(\a1/k1a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [30]),
        .Q(\a1/k1a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [31]),
        .Q(\a1/k1a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [3]),
        .Q(\a1/k1a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [4]),
        .Q(\a1/k1a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [5]),
        .Q(\a1/k1a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [6]),
        .Q(\a1/k1a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [7]),
        .Q(\a1/k1a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [8]),
        .Q(\a1/k1a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k1a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v1 [9]),
        .Q(\a1/k1a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [0]),
        .Q(\a1/k2a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [10]),
        .Q(\a1/k2a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [11]),
        .Q(\a1/k2a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [12]),
        .Q(\a1/k2a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [13]),
        .Q(\a1/k2a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [14]),
        .Q(\a1/k2a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [15]),
        .Q(\a1/k2a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [16]),
        .Q(\a1/k2a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [17]),
        .Q(\a1/k2a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [18]),
        .Q(\a1/k2a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [19]),
        .Q(\a1/k2a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [1]),
        .Q(\a1/k2a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [20]),
        .Q(\a1/k2a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [21]),
        .Q(\a1/k2a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [22]),
        .Q(\a1/k2a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [23]),
        .Q(\a1/k2a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [24]),
        .Q(\a1/k2a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [25]),
        .Q(\a1/k2a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [26]),
        .Q(\a1/k2a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [27]),
        .Q(\a1/k2a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [28]),
        .Q(\a1/k2a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [29]),
        .Q(\a1/k2a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [2]),
        .Q(\a1/k2a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [30]),
        .Q(\a1/k2a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [31]),
        .Q(\a1/k2a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [3]),
        .Q(\a1/k2a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [4]),
        .Q(\a1/k2a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [5]),
        .Q(\a1/k2a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [6]),
        .Q(\a1/k2a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [7]),
        .Q(\a1/k2a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [8]),
        .Q(\a1/k2a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k2a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v2 [9]),
        .Q(\a1/k2a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [0]),
        .Q(\a1/k3a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [10]),
        .Q(\a1/k3a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [11]),
        .Q(\a1/k3a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [12]),
        .Q(\a1/k3a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [13]),
        .Q(\a1/k3a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [14]),
        .Q(\a1/k3a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [15]),
        .Q(\a1/k3a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [16]),
        .Q(\a1/k3a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [17]),
        .Q(\a1/k3a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [18]),
        .Q(\a1/k3a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [19]),
        .Q(\a1/k3a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [1]),
        .Q(\a1/k3a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [20]),
        .Q(\a1/k3a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [21]),
        .Q(\a1/k3a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [22]),
        .Q(\a1/k3a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [23]),
        .Q(\a1/k3a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [24]),
        .Q(\a1/k3a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [25]),
        .Q(\a1/k3a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [26]),
        .Q(\a1/k3a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [27]),
        .Q(\a1/k3a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [28]),
        .Q(\a1/k3a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [29]),
        .Q(\a1/k3a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [2]),
        .Q(\a1/k3a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [30]),
        .Q(\a1/k3a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [31]),
        .Q(\a1/k3a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [3]),
        .Q(\a1/k3a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [4]),
        .Q(\a1/k3a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [5]),
        .Q(\a1/k3a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [6]),
        .Q(\a1/k3a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [7]),
        .Q(\a1/k3a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [8]),
        .Q(\a1/k3a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/k3a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a1/v3 [9]),
        .Q(\a1/k3a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[0]),
        .Q(k1[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[100] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[100]),
        .Q(k1[100]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[101] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[101]),
        .Q(k1[101]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[102] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[102]),
        .Q(k1[102]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[103] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[103]),
        .Q(k1[103]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[104] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[104]),
        .Q(k1[104]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[105] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[105]),
        .Q(k1[105]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[106] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[106]),
        .Q(k1[106]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[107] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[107]),
        .Q(k1[107]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[108] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[108]),
        .Q(k1[108]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[109] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[109]),
        .Q(k1[109]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[10]),
        .Q(k1[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[110] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[110]),
        .Q(k1[110]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[111] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[111]),
        .Q(k1[111]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[112] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[112]),
        .Q(k1[112]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[113] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[113]),
        .Q(k1[113]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[114] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[114]),
        .Q(k1[114]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[115] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[115]),
        .Q(k1[115]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[116] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[116]),
        .Q(k1[116]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[117] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[117]),
        .Q(k1[117]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[118] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[118]),
        .Q(k1[118]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[119] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[119]),
        .Q(k1[119]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[11]),
        .Q(k1[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[120] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[120]),
        .Q(k1[120]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[121] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[121]),
        .Q(k1[121]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[122] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[122]),
        .Q(k1[122]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[123] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[123]),
        .Q(k1[123]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[124] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[124]),
        .Q(k1[124]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[125] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[125]),
        .Q(k1[125]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[126] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[126]),
        .Q(k1[126]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[127] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[127]),
        .Q(k1[127]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[12]),
        .Q(k1[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[13]),
        .Q(k1[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[14]),
        .Q(k1[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[15]),
        .Q(k1[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[16]),
        .Q(k1[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[17]),
        .Q(k1[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[18]),
        .Q(k1[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[19]),
        .Q(k1[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[1]),
        .Q(k1[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[20]),
        .Q(k1[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[21]),
        .Q(k1[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[22]),
        .Q(k1[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[23]),
        .Q(k1[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[24]),
        .Q(k1[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[25]),
        .Q(k1[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[26]),
        .Q(k1[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[27]),
        .Q(k1[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[28]),
        .Q(k1[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[29]),
        .Q(k1[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[2]),
        .Q(k1[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[30]),
        .Q(k1[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[31]),
        .Q(k1[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[32]),
        .Q(k1[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[33]),
        .Q(k1[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[34]),
        .Q(k1[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[35]),
        .Q(k1[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[36]),
        .Q(k1[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[37]),
        .Q(k1[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[38]),
        .Q(k1[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[39]),
        .Q(k1[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[3]),
        .Q(k1[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[40]),
        .Q(k1[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[41]),
        .Q(k1[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[42]),
        .Q(k1[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[43]),
        .Q(k1[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[44]),
        .Q(k1[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[45]),
        .Q(k1[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[46]),
        .Q(k1[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[47]),
        .Q(k1[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[48]),
        .Q(k1[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[49]),
        .Q(k1[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[4]),
        .Q(k1[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[50]),
        .Q(k1[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[51]),
        .Q(k1[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[52]),
        .Q(k1[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[53]),
        .Q(k1[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[54]),
        .Q(k1[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[55]),
        .Q(k1[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[56]),
        .Q(k1[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[57]),
        .Q(k1[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[58]),
        .Q(k1[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[59]),
        .Q(k1[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[5]),
        .Q(k1[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[60]),
        .Q(k1[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[61]),
        .Q(k1[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[62]),
        .Q(k1[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[63]),
        .Q(k1[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[64] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[64]),
        .Q(k1[64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[65] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[65]),
        .Q(k1[65]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[66] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[66]),
        .Q(k1[66]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[67] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[67]),
        .Q(k1[67]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[68] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[68]),
        .Q(k1[68]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[69] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[69]),
        .Q(k1[69]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[6]),
        .Q(k1[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[70] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[70]),
        .Q(k1[70]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[71] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[71]),
        .Q(k1[71]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[72] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[72]),
        .Q(k1[72]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[73] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[73]),
        .Q(k1[73]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[74] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[74]),
        .Q(k1[74]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[75] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[75]),
        .Q(k1[75]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[76] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[76]),
        .Q(k1[76]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[77] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[77]),
        .Q(k1[77]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[78] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[78]),
        .Q(k1[78]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[79] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[79]),
        .Q(k1[79]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[7]),
        .Q(k1[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[80] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[80]),
        .Q(k1[80]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[81] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[81]),
        .Q(k1[81]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[82] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[82]),
        .Q(k1[82]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[83] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[83]),
        .Q(k1[83]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[84] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[84]),
        .Q(k1[84]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[85] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[85]),
        .Q(k1[85]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[86] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[86]),
        .Q(k1[86]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[87] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[87]),
        .Q(k1[87]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[88] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[88]),
        .Q(k1[88]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[89] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[89]),
        .Q(k1[89]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[8]),
        .Q(k1[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[90] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[90]),
        .Q(k1[90]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[91] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[91]),
        .Q(k1[91]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[92] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[92]),
        .Q(k1[92]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[93] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[93]),
        .Q(k1[93]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[94] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[94]),
        .Q(k1[94]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[95] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[95]),
        .Q(k1[95]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[96] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[96]),
        .Q(k1[96]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[97] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[97]),
        .Q(k1[97]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[98] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[98]),
        .Q(k1[98]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[99] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[99]),
        .Q(k1[99]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a1/out_1_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k0b[9]),
        .Q(k1[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_0/S_1/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \a10/S4_0/S_1/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,k9[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,k9[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\a10/S4_0/S_1/out_reg_n_0 ,\a10/S4_0/S_1/out_reg_n_1 ,\a10/S4_0/S_1/out_reg_n_2 ,\a10/S4_0/S_1/out_reg_n_3 ,\a10/S4_0/S_1/out_reg_n_4 ,\a10/S4_0/S_1/out_reg_n_5 ,\a10/S4_0/S_1/out_reg_n_6 ,\a10/S4_0/S_1/out_reg_n_7 ,\a10/k4a [23:16]}),
        .DOBDO({\a10/S4_0/S_1/out_reg_n_16 ,\a10/S4_0/S_1/out_reg_n_17 ,\a10/S4_0/S_1/out_reg_n_18 ,\a10/S4_0/S_1/out_reg_n_19 ,\a10/S4_0/S_1/out_reg_n_20 ,\a10/S4_0/S_1/out_reg_n_21 ,\a10/S4_0/S_1/out_reg_n_22 ,\a10/S4_0/S_1/out_reg_n_23 ,\a10/k4a [31:24]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_0/S_3/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \a10/S4_0/S_3/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,k9[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,k9[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\a10/S4_0/S_3/out_reg_n_0 ,\a10/S4_0/S_3/out_reg_n_1 ,\a10/S4_0/S_3/out_reg_n_2 ,\a10/S4_0/S_3/out_reg_n_3 ,\a10/S4_0/S_3/out_reg_n_4 ,\a10/S4_0/S_3/out_reg_n_5 ,\a10/S4_0/S_3/out_reg_n_6 ,\a10/S4_0/S_3/out_reg_n_7 ,\a10/k4a [7:0]}),
        .DOBDO({\a10/S4_0/S_3/out_reg_n_16 ,\a10/S4_0/S_3/out_reg_n_17 ,\a10/S4_0/S_3/out_reg_n_18 ,\a10/S4_0/S_3/out_reg_n_19 ,\a10/S4_0/S_3/out_reg_n_20 ,\a10/S4_0/S_3/out_reg_n_21 ,\a10/S4_0/S_3/out_reg_n_22 ,\a10/S4_0/S_3/out_reg_n_23 ,\a10/k4a [15:8]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[96]),
        .Q(\a10/k0a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[106]),
        .Q(\a10/k0a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[107]),
        .Q(\a10/k0a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[108]),
        .Q(\a10/k0a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[109]),
        .Q(\a10/k0a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[110]),
        .Q(\a10/k0a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[111]),
        .Q(\a10/k0a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[112]),
        .Q(\a10/k0a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[113]),
        .Q(\a10/k0a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[114]),
        .Q(\a10/k0a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[115]),
        .Q(\a10/k0a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[97]),
        .Q(\a10/k0a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[116]),
        .Q(\a10/k0a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[117]),
        .Q(\a10/k0a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[118]),
        .Q(\a10/k0a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[119]),
        .Q(\a10/k0a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[120]),
        .Q(\a10/k0a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v0 [25]),
        .Q(\a10/k0a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v0 [26]),
        .Q(\a10/k0a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[123]),
        .Q(\a10/k0a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v0 [28]),
        .Q(\a10/k0a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v0 [29]),
        .Q(\a10/k0a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[98]),
        .Q(\a10/k0a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[126]),
        .Q(\a10/k0a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[127]),
        .Q(\a10/k0a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[99]),
        .Q(\a10/k0a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[100]),
        .Q(\a10/k0a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[101]),
        .Q(\a10/k0a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[102]),
        .Q(\a10/k0a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[103]),
        .Q(\a10/k0a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[104]),
        .Q(\a10/k0a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k0a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k9[105]),
        .Q(\a10/k0a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [0]),
        .Q(\a10/k1a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [10]),
        .Q(\a10/k1a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [11]),
        .Q(\a10/k1a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [12]),
        .Q(\a10/k1a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [13]),
        .Q(\a10/k1a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [14]),
        .Q(\a10/k1a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [15]),
        .Q(\a10/k1a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [16]),
        .Q(\a10/k1a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [17]),
        .Q(\a10/k1a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [18]),
        .Q(\a10/k1a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [19]),
        .Q(\a10/k1a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [1]),
        .Q(\a10/k1a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [20]),
        .Q(\a10/k1a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [21]),
        .Q(\a10/k1a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [22]),
        .Q(\a10/k1a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [23]),
        .Q(\a10/k1a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [24]),
        .Q(\a10/k1a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\k1a[25]_i_1__8_n_0 ),
        .Q(\a10/k1a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\k1a[26]_i_1__8_n_0 ),
        .Q(\a10/k1a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [27]),
        .Q(\a10/k1a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\k1a[28]_i_1__8_n_0 ),
        .Q(\a10/k1a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\k1a[29]_i_1__8_n_0 ),
        .Q(\a10/k1a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [2]),
        .Q(\a10/k1a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [30]),
        .Q(\a10/k1a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [31]),
        .Q(\a10/k1a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [3]),
        .Q(\a10/k1a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [4]),
        .Q(\a10/k1a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [5]),
        .Q(\a10/k1a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [6]),
        .Q(\a10/k1a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [7]),
        .Q(\a10/k1a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [8]),
        .Q(\a10/k1a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k1a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v1 [9]),
        .Q(\a10/k1a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [0]),
        .Q(\a10/k2a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [10]),
        .Q(\a10/k2a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [11]),
        .Q(\a10/k2a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [12]),
        .Q(\a10/k2a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [13]),
        .Q(\a10/k2a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [14]),
        .Q(\a10/k2a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [15]),
        .Q(\a10/k2a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [16]),
        .Q(\a10/k2a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [17]),
        .Q(\a10/k2a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [18]),
        .Q(\a10/k2a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [19]),
        .Q(\a10/k2a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [1]),
        .Q(\a10/k2a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [20]),
        .Q(\a10/k2a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [21]),
        .Q(\a10/k2a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [22]),
        .Q(\a10/k2a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [23]),
        .Q(\a10/k2a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [24]),
        .Q(\a10/k2a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [25]),
        .Q(\a10/k2a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [26]),
        .Q(\a10/k2a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [27]),
        .Q(\a10/k2a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [28]),
        .Q(\a10/k2a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [29]),
        .Q(\a10/k2a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [2]),
        .Q(\a10/k2a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [30]),
        .Q(\a10/k2a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [31]),
        .Q(\a10/k2a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [3]),
        .Q(\a10/k2a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [4]),
        .Q(\a10/k2a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [5]),
        .Q(\a10/k2a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [6]),
        .Q(\a10/k2a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [7]),
        .Q(\a10/k2a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [8]),
        .Q(\a10/k2a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k2a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v2 [9]),
        .Q(\a10/k2a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [0]),
        .Q(\a10/k3a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [10]),
        .Q(\a10/k3a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [11]),
        .Q(\a10/k3a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [12]),
        .Q(\a10/k3a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [13]),
        .Q(\a10/k3a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [14]),
        .Q(\a10/k3a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [15]),
        .Q(\a10/k3a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [16]),
        .Q(\a10/k3a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [17]),
        .Q(\a10/k3a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [18]),
        .Q(\a10/k3a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [19]),
        .Q(\a10/k3a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [1]),
        .Q(\a10/k3a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [20]),
        .Q(\a10/k3a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [21]),
        .Q(\a10/k3a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [22]),
        .Q(\a10/k3a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [23]),
        .Q(\a10/k3a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [24]),
        .Q(\a10/k3a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [25]),
        .Q(\a10/k3a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [26]),
        .Q(\a10/k3a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [27]),
        .Q(\a10/k3a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [28]),
        .Q(\a10/k3a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [29]),
        .Q(\a10/k3a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [2]),
        .Q(\a10/k3a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [30]),
        .Q(\a10/k3a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [31]),
        .Q(\a10/k3a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [3]),
        .Q(\a10/k3a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [4]),
        .Q(\a10/k3a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [5]),
        .Q(\a10/k3a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [6]),
        .Q(\a10/k3a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [7]),
        .Q(\a10/k3a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [8]),
        .Q(\a10/k3a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a10/k3a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a10/v3 [9]),
        .Q(\a10/k3a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_0/S_1/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \a2/S4_0/S_1/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,k1[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,k1[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\a2/S4_0/S_1/out_reg_n_0 ,\a2/S4_0/S_1/out_reg_n_1 ,\a2/S4_0/S_1/out_reg_n_2 ,\a2/S4_0/S_1/out_reg_n_3 ,\a2/S4_0/S_1/out_reg_n_4 ,\a2/S4_0/S_1/out_reg_n_5 ,\a2/S4_0/S_1/out_reg_n_6 ,\a2/S4_0/S_1/out_reg_n_7 ,\a2/k4a [23:16]}),
        .DOBDO({\a2/S4_0/S_1/out_reg_n_16 ,\a2/S4_0/S_1/out_reg_n_17 ,\a2/S4_0/S_1/out_reg_n_18 ,\a2/S4_0/S_1/out_reg_n_19 ,\a2/S4_0/S_1/out_reg_n_20 ,\a2/S4_0/S_1/out_reg_n_21 ,\a2/S4_0/S_1/out_reg_n_22 ,\a2/S4_0/S_1/out_reg_n_23 ,\a2/k4a [31:24]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_0/S_3/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \a2/S4_0/S_3/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,k1[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,k1[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\a2/S4_0/S_3/out_reg_n_0 ,\a2/S4_0/S_3/out_reg_n_1 ,\a2/S4_0/S_3/out_reg_n_2 ,\a2/S4_0/S_3/out_reg_n_3 ,\a2/S4_0/S_3/out_reg_n_4 ,\a2/S4_0/S_3/out_reg_n_5 ,\a2/S4_0/S_3/out_reg_n_6 ,\a2/S4_0/S_3/out_reg_n_7 ,\a2/k4a [7:0]}),
        .DOBDO({\a2/S4_0/S_3/out_reg_n_16 ,\a2/S4_0/S_3/out_reg_n_17 ,\a2/S4_0/S_3/out_reg_n_18 ,\a2/S4_0/S_3/out_reg_n_19 ,\a2/S4_0/S_3/out_reg_n_20 ,\a2/S4_0/S_3/out_reg_n_21 ,\a2/S4_0/S_3/out_reg_n_22 ,\a2/S4_0/S_3/out_reg_n_23 ,\a2/k4a [15:8]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[96]),
        .Q(\a2/k0a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[106]),
        .Q(\a2/k0a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[107]),
        .Q(\a2/k0a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[108]),
        .Q(\a2/k0a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[109]),
        .Q(\a2/k0a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[110]),
        .Q(\a2/k0a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[111]),
        .Q(\a2/k0a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[112]),
        .Q(\a2/k0a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[113]),
        .Q(\a2/k0a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[114]),
        .Q(\a2/k0a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[115]),
        .Q(\a2/k0a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[97]),
        .Q(\a2/k0a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[116]),
        .Q(\a2/k0a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[117]),
        .Q(\a2/k0a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[118]),
        .Q(\a2/k0a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[119]),
        .Q(\a2/k0a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[120]),
        .Q(\a2/k0a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v0 ),
        .Q(\a2/k0a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[122]),
        .Q(\a2/k0a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[123]),
        .Q(\a2/k0a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[124]),
        .Q(\a2/k0a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[125]),
        .Q(\a2/k0a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[98]),
        .Q(\a2/k0a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[126]),
        .Q(\a2/k0a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[127]),
        .Q(\a2/k0a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[99]),
        .Q(\a2/k0a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[100]),
        .Q(\a2/k0a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[101]),
        .Q(\a2/k0a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[102]),
        .Q(\a2/k0a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[103]),
        .Q(\a2/k0a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[104]),
        .Q(\a2/k0a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k0a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1[105]),
        .Q(\a2/k0a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [0]),
        .Q(\a2/k1a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [10]),
        .Q(\a2/k1a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [11]),
        .Q(\a2/k1a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [12]),
        .Q(\a2/k1a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [13]),
        .Q(\a2/k1a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [14]),
        .Q(\a2/k1a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [15]),
        .Q(\a2/k1a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [16]),
        .Q(\a2/k1a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [17]),
        .Q(\a2/k1a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [18]),
        .Q(\a2/k1a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [19]),
        .Q(\a2/k1a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [1]),
        .Q(\a2/k1a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [20]),
        .Q(\a2/k1a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [21]),
        .Q(\a2/k1a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [22]),
        .Q(\a2/k1a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [23]),
        .Q(\a2/k1a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [24]),
        .Q(\a2/k1a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\k1a[25]_i_1__0_n_0 ),
        .Q(\a2/k1a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [26]),
        .Q(\a2/k1a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [27]),
        .Q(\a2/k1a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [28]),
        .Q(\a2/k1a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [29]),
        .Q(\a2/k1a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [2]),
        .Q(\a2/k1a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [30]),
        .Q(\a2/k1a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [31]),
        .Q(\a2/k1a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [3]),
        .Q(\a2/k1a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [4]),
        .Q(\a2/k1a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [5]),
        .Q(\a2/k1a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [6]),
        .Q(\a2/k1a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [7]),
        .Q(\a2/k1a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [8]),
        .Q(\a2/k1a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k1a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v1 [9]),
        .Q(\a2/k1a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [0]),
        .Q(\a2/k2a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [10]),
        .Q(\a2/k2a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [11]),
        .Q(\a2/k2a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [12]),
        .Q(\a2/k2a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [13]),
        .Q(\a2/k2a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [14]),
        .Q(\a2/k2a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [15]),
        .Q(\a2/k2a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [16]),
        .Q(\a2/k2a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [17]),
        .Q(\a2/k2a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [18]),
        .Q(\a2/k2a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [19]),
        .Q(\a2/k2a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [1]),
        .Q(\a2/k2a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [20]),
        .Q(\a2/k2a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [21]),
        .Q(\a2/k2a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [22]),
        .Q(\a2/k2a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [23]),
        .Q(\a2/k2a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [24]),
        .Q(\a2/k2a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [25]),
        .Q(\a2/k2a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [26]),
        .Q(\a2/k2a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [27]),
        .Q(\a2/k2a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [28]),
        .Q(\a2/k2a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [29]),
        .Q(\a2/k2a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [2]),
        .Q(\a2/k2a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [30]),
        .Q(\a2/k2a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [31]),
        .Q(\a2/k2a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [3]),
        .Q(\a2/k2a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [4]),
        .Q(\a2/k2a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [5]),
        .Q(\a2/k2a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [6]),
        .Q(\a2/k2a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [7]),
        .Q(\a2/k2a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [8]),
        .Q(\a2/k2a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k2a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v2 [9]),
        .Q(\a2/k2a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [0]),
        .Q(\a2/k3a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [10]),
        .Q(\a2/k3a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [11]),
        .Q(\a2/k3a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [12]),
        .Q(\a2/k3a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [13]),
        .Q(\a2/k3a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [14]),
        .Q(\a2/k3a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [15]),
        .Q(\a2/k3a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [16]),
        .Q(\a2/k3a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [17]),
        .Q(\a2/k3a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [18]),
        .Q(\a2/k3a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [19]),
        .Q(\a2/k3a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [1]),
        .Q(\a2/k3a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [20]),
        .Q(\a2/k3a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [21]),
        .Q(\a2/k3a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [22]),
        .Q(\a2/k3a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [23]),
        .Q(\a2/k3a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [24]),
        .Q(\a2/k3a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [25]),
        .Q(\a2/k3a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [26]),
        .Q(\a2/k3a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [27]),
        .Q(\a2/k3a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [28]),
        .Q(\a2/k3a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [29]),
        .Q(\a2/k3a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [2]),
        .Q(\a2/k3a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [30]),
        .Q(\a2/k3a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [31]),
        .Q(\a2/k3a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [3]),
        .Q(\a2/k3a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [4]),
        .Q(\a2/k3a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [5]),
        .Q(\a2/k3a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [6]),
        .Q(\a2/k3a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [7]),
        .Q(\a2/k3a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [8]),
        .Q(\a2/k3a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/k3a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a2/v3 [9]),
        .Q(\a2/k3a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[0]),
        .Q(k2[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[100] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[100]),
        .Q(k2[100]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[101] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[101]),
        .Q(k2[101]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[102] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[102]),
        .Q(k2[102]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[103] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[103]),
        .Q(k2[103]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[104] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[104]),
        .Q(k2[104]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[105] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[105]),
        .Q(k2[105]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[106] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[106]),
        .Q(k2[106]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[107] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[107]),
        .Q(k2[107]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[108] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[108]),
        .Q(k2[108]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[109] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[109]),
        .Q(k2[109]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[10]),
        .Q(k2[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[110] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[110]),
        .Q(k2[110]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[111] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[111]),
        .Q(k2[111]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[112] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[112]),
        .Q(k2[112]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[113] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[113]),
        .Q(k2[113]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[114] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[114]),
        .Q(k2[114]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[115] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[115]),
        .Q(k2[115]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[116] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[116]),
        .Q(k2[116]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[117] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[117]),
        .Q(k2[117]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[118] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[118]),
        .Q(k2[118]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[119] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[119]),
        .Q(k2[119]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[11]),
        .Q(k2[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[120] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[120]),
        .Q(k2[120]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[121] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[121]),
        .Q(k2[121]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[122] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[122]),
        .Q(k2[122]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[123] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[123]),
        .Q(k2[123]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[124] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[124]),
        .Q(k2[124]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[125] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[125]),
        .Q(k2[125]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[126] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[126]),
        .Q(k2[126]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[127] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[127]),
        .Q(k2[127]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[12]),
        .Q(k2[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[13]),
        .Q(k2[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[14]),
        .Q(k2[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[15]),
        .Q(k2[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[16]),
        .Q(k2[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[17]),
        .Q(k2[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[18]),
        .Q(k2[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[19]),
        .Q(k2[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[1]),
        .Q(k2[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[20]),
        .Q(k2[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[21]),
        .Q(k2[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[22]),
        .Q(k2[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[23]),
        .Q(k2[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[24]),
        .Q(k2[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[25]),
        .Q(k2[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[26]),
        .Q(k2[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[27]),
        .Q(k2[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[28]),
        .Q(k2[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[29]),
        .Q(k2[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[2]),
        .Q(k2[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[30]),
        .Q(k2[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[31]),
        .Q(k2[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[32]),
        .Q(k2[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[33]),
        .Q(k2[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[34]),
        .Q(k2[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[35]),
        .Q(k2[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[36]),
        .Q(k2[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[37]),
        .Q(k2[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[38]),
        .Q(k2[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[39]),
        .Q(k2[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[3]),
        .Q(k2[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[40]),
        .Q(k2[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[41]),
        .Q(k2[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[42]),
        .Q(k2[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[43]),
        .Q(k2[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[44]),
        .Q(k2[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[45]),
        .Q(k2[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[46]),
        .Q(k2[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[47]),
        .Q(k2[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[48]),
        .Q(k2[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[49]),
        .Q(k2[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[4]),
        .Q(k2[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[50]),
        .Q(k2[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[51]),
        .Q(k2[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[52]),
        .Q(k2[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[53]),
        .Q(k2[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[54]),
        .Q(k2[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[55]),
        .Q(k2[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[56]),
        .Q(k2[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[57]),
        .Q(k2[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[58]),
        .Q(k2[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[59]),
        .Q(k2[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[5]),
        .Q(k2[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[60]),
        .Q(k2[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[61]),
        .Q(k2[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[62]),
        .Q(k2[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[63]),
        .Q(k2[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[64] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[64]),
        .Q(k2[64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[65] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[65]),
        .Q(k2[65]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[66] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[66]),
        .Q(k2[66]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[67] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[67]),
        .Q(k2[67]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[68] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[68]),
        .Q(k2[68]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[69] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[69]),
        .Q(k2[69]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[6]),
        .Q(k2[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[70] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[70]),
        .Q(k2[70]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[71] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[71]),
        .Q(k2[71]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[72] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[72]),
        .Q(k2[72]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[73] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[73]),
        .Q(k2[73]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[74] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[74]),
        .Q(k2[74]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[75] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[75]),
        .Q(k2[75]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[76] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[76]),
        .Q(k2[76]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[77] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[77]),
        .Q(k2[77]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[78] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[78]),
        .Q(k2[78]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[79] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[79]),
        .Q(k2[79]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[7]),
        .Q(k2[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[80] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[80]),
        .Q(k2[80]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[81] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[81]),
        .Q(k2[81]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[82] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[82]),
        .Q(k2[82]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[83] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[83]),
        .Q(k2[83]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[84] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[84]),
        .Q(k2[84]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[85] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[85]),
        .Q(k2[85]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[86] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[86]),
        .Q(k2[86]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[87] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[87]),
        .Q(k2[87]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[88] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[88]),
        .Q(k2[88]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[89] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[89]),
        .Q(k2[89]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[8]),
        .Q(k2[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[90] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[90]),
        .Q(k2[90]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[91] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[91]),
        .Q(k2[91]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[92] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[92]),
        .Q(k2[92]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[93] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[93]),
        .Q(k2[93]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[94] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[94]),
        .Q(k2[94]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[95] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[95]),
        .Q(k2[95]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[96] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[96]),
        .Q(k2[96]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[97] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[97]),
        .Q(k2[97]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[98] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[98]),
        .Q(k2[98]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[99] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[99]),
        .Q(k2[99]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a2/out_1_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1b[9]),
        .Q(k2[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_0/S_1/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \a3/S4_0/S_1/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,k2[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,k2[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\a3/S4_0/S_1/out_reg_n_0 ,\a3/S4_0/S_1/out_reg_n_1 ,\a3/S4_0/S_1/out_reg_n_2 ,\a3/S4_0/S_1/out_reg_n_3 ,\a3/S4_0/S_1/out_reg_n_4 ,\a3/S4_0/S_1/out_reg_n_5 ,\a3/S4_0/S_1/out_reg_n_6 ,\a3/S4_0/S_1/out_reg_n_7 ,\a3/k4a [23:16]}),
        .DOBDO({\a3/S4_0/S_1/out_reg_n_16 ,\a3/S4_0/S_1/out_reg_n_17 ,\a3/S4_0/S_1/out_reg_n_18 ,\a3/S4_0/S_1/out_reg_n_19 ,\a3/S4_0/S_1/out_reg_n_20 ,\a3/S4_0/S_1/out_reg_n_21 ,\a3/S4_0/S_1/out_reg_n_22 ,\a3/S4_0/S_1/out_reg_n_23 ,\a3/k4a [31:24]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_0/S_3/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \a3/S4_0/S_3/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,k2[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,k2[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\a3/S4_0/S_3/out_reg_n_0 ,\a3/S4_0/S_3/out_reg_n_1 ,\a3/S4_0/S_3/out_reg_n_2 ,\a3/S4_0/S_3/out_reg_n_3 ,\a3/S4_0/S_3/out_reg_n_4 ,\a3/S4_0/S_3/out_reg_n_5 ,\a3/S4_0/S_3/out_reg_n_6 ,\a3/S4_0/S_3/out_reg_n_7 ,\a3/k4a [7:0]}),
        .DOBDO({\a3/S4_0/S_3/out_reg_n_16 ,\a3/S4_0/S_3/out_reg_n_17 ,\a3/S4_0/S_3/out_reg_n_18 ,\a3/S4_0/S_3/out_reg_n_19 ,\a3/S4_0/S_3/out_reg_n_20 ,\a3/S4_0/S_3/out_reg_n_21 ,\a3/S4_0/S_3/out_reg_n_22 ,\a3/S4_0/S_3/out_reg_n_23 ,\a3/k4a [15:8]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[96]),
        .Q(\a3/k0a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[106]),
        .Q(\a3/k0a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[107]),
        .Q(\a3/k0a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[108]),
        .Q(\a3/k0a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[109]),
        .Q(\a3/k0a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[110]),
        .Q(\a3/k0a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[111]),
        .Q(\a3/k0a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[112]),
        .Q(\a3/k0a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[113]),
        .Q(\a3/k0a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[114]),
        .Q(\a3/k0a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[115]),
        .Q(\a3/k0a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[97]),
        .Q(\a3/k0a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[116]),
        .Q(\a3/k0a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[117]),
        .Q(\a3/k0a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[118]),
        .Q(\a3/k0a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[119]),
        .Q(\a3/k0a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[120]),
        .Q(\a3/k0a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[121]),
        .Q(\a3/k0a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v0 ),
        .Q(\a3/k0a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[123]),
        .Q(\a3/k0a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[124]),
        .Q(\a3/k0a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[125]),
        .Q(\a3/k0a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[98]),
        .Q(\a3/k0a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[126]),
        .Q(\a3/k0a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[127]),
        .Q(\a3/k0a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[99]),
        .Q(\a3/k0a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[100]),
        .Q(\a3/k0a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[101]),
        .Q(\a3/k0a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[102]),
        .Q(\a3/k0a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[103]),
        .Q(\a3/k0a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[104]),
        .Q(\a3/k0a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k0a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2[105]),
        .Q(\a3/k0a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [0]),
        .Q(\a3/k1a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [10]),
        .Q(\a3/k1a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [11]),
        .Q(\a3/k1a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [12]),
        .Q(\a3/k1a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [13]),
        .Q(\a3/k1a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [14]),
        .Q(\a3/k1a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [15]),
        .Q(\a3/k1a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [16]),
        .Q(\a3/k1a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [17]),
        .Q(\a3/k1a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [18]),
        .Q(\a3/k1a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [19]),
        .Q(\a3/k1a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [1]),
        .Q(\a3/k1a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [20]),
        .Q(\a3/k1a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [21]),
        .Q(\a3/k1a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [22]),
        .Q(\a3/k1a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [23]),
        .Q(\a3/k1a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [24]),
        .Q(\a3/k1a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [25]),
        .Q(\a3/k1a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\k1a[26]_i_1__1_n_0 ),
        .Q(\a3/k1a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [27]),
        .Q(\a3/k1a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [28]),
        .Q(\a3/k1a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [29]),
        .Q(\a3/k1a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [2]),
        .Q(\a3/k1a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [30]),
        .Q(\a3/k1a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [31]),
        .Q(\a3/k1a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [3]),
        .Q(\a3/k1a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [4]),
        .Q(\a3/k1a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [5]),
        .Q(\a3/k1a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [6]),
        .Q(\a3/k1a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [7]),
        .Q(\a3/k1a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [8]),
        .Q(\a3/k1a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k1a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v1 [9]),
        .Q(\a3/k1a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [0]),
        .Q(\a3/k2a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [10]),
        .Q(\a3/k2a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [11]),
        .Q(\a3/k2a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [12]),
        .Q(\a3/k2a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [13]),
        .Q(\a3/k2a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [14]),
        .Q(\a3/k2a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [15]),
        .Q(\a3/k2a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [16]),
        .Q(\a3/k2a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [17]),
        .Q(\a3/k2a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [18]),
        .Q(\a3/k2a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [19]),
        .Q(\a3/k2a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [1]),
        .Q(\a3/k2a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [20]),
        .Q(\a3/k2a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [21]),
        .Q(\a3/k2a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [22]),
        .Q(\a3/k2a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [23]),
        .Q(\a3/k2a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [24]),
        .Q(\a3/k2a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [25]),
        .Q(\a3/k2a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [26]),
        .Q(\a3/k2a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [27]),
        .Q(\a3/k2a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [28]),
        .Q(\a3/k2a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [29]),
        .Q(\a3/k2a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [2]),
        .Q(\a3/k2a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [30]),
        .Q(\a3/k2a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [31]),
        .Q(\a3/k2a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [3]),
        .Q(\a3/k2a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [4]),
        .Q(\a3/k2a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [5]),
        .Q(\a3/k2a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [6]),
        .Q(\a3/k2a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [7]),
        .Q(\a3/k2a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [8]),
        .Q(\a3/k2a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k2a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v2 [9]),
        .Q(\a3/k2a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [0]),
        .Q(\a3/k3a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [10]),
        .Q(\a3/k3a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [11]),
        .Q(\a3/k3a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [12]),
        .Q(\a3/k3a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [13]),
        .Q(\a3/k3a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [14]),
        .Q(\a3/k3a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [15]),
        .Q(\a3/k3a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [16]),
        .Q(\a3/k3a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [17]),
        .Q(\a3/k3a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [18]),
        .Q(\a3/k3a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [19]),
        .Q(\a3/k3a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [1]),
        .Q(\a3/k3a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [20]),
        .Q(\a3/k3a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [21]),
        .Q(\a3/k3a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [22]),
        .Q(\a3/k3a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [23]),
        .Q(\a3/k3a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [24]),
        .Q(\a3/k3a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [25]),
        .Q(\a3/k3a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [26]),
        .Q(\a3/k3a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [27]),
        .Q(\a3/k3a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [28]),
        .Q(\a3/k3a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [29]),
        .Q(\a3/k3a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [2]),
        .Q(\a3/k3a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [30]),
        .Q(\a3/k3a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [31]),
        .Q(\a3/k3a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [3]),
        .Q(\a3/k3a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [4]),
        .Q(\a3/k3a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [5]),
        .Q(\a3/k3a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [6]),
        .Q(\a3/k3a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [7]),
        .Q(\a3/k3a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [8]),
        .Q(\a3/k3a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/k3a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a3/v3 [9]),
        .Q(\a3/k3a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[0]),
        .Q(k3[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[100] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[100]),
        .Q(k3[100]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[101] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[101]),
        .Q(k3[101]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[102] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[102]),
        .Q(k3[102]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[103] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[103]),
        .Q(k3[103]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[104] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[104]),
        .Q(k3[104]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[105] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[105]),
        .Q(k3[105]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[106] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[106]),
        .Q(k3[106]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[107] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[107]),
        .Q(k3[107]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[108] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[108]),
        .Q(k3[108]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[109] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[109]),
        .Q(k3[109]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[10]),
        .Q(k3[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[110] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[110]),
        .Q(k3[110]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[111] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[111]),
        .Q(k3[111]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[112] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[112]),
        .Q(k3[112]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[113] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[113]),
        .Q(k3[113]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[114] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[114]),
        .Q(k3[114]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[115] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[115]),
        .Q(k3[115]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[116] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[116]),
        .Q(k3[116]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[117] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[117]),
        .Q(k3[117]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[118] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[118]),
        .Q(k3[118]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[119] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[119]),
        .Q(k3[119]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[11]),
        .Q(k3[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[120] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[120]),
        .Q(k3[120]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[121] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[121]),
        .Q(k3[121]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[122] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[122]),
        .Q(k3[122]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[123] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[123]),
        .Q(k3[123]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[124] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[124]),
        .Q(k3[124]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[125] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[125]),
        .Q(k3[125]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[126] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[126]),
        .Q(k3[126]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[127] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[127]),
        .Q(k3[127]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[12]),
        .Q(k3[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[13]),
        .Q(k3[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[14]),
        .Q(k3[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[15]),
        .Q(k3[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[16]),
        .Q(k3[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[17]),
        .Q(k3[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[18]),
        .Q(k3[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[19]),
        .Q(k3[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[1]),
        .Q(k3[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[20]),
        .Q(k3[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[21]),
        .Q(k3[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[22]),
        .Q(k3[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[23]),
        .Q(k3[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[24]),
        .Q(k3[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[25]),
        .Q(k3[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[26]),
        .Q(k3[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[27]),
        .Q(k3[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[28]),
        .Q(k3[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[29]),
        .Q(k3[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[2]),
        .Q(k3[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[30]),
        .Q(k3[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[31]),
        .Q(k3[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[32]),
        .Q(k3[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[33]),
        .Q(k3[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[34]),
        .Q(k3[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[35]),
        .Q(k3[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[36]),
        .Q(k3[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[37]),
        .Q(k3[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[38]),
        .Q(k3[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[39]),
        .Q(k3[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[3]),
        .Q(k3[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[40]),
        .Q(k3[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[41]),
        .Q(k3[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[42]),
        .Q(k3[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[43]),
        .Q(k3[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[44]),
        .Q(k3[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[45]),
        .Q(k3[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[46]),
        .Q(k3[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[47]),
        .Q(k3[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[48]),
        .Q(k3[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[49]),
        .Q(k3[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[4]),
        .Q(k3[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[50]),
        .Q(k3[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[51]),
        .Q(k3[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[52]),
        .Q(k3[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[53]),
        .Q(k3[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[54]),
        .Q(k3[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[55]),
        .Q(k3[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[56]),
        .Q(k3[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[57]),
        .Q(k3[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[58]),
        .Q(k3[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[59]),
        .Q(k3[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[5]),
        .Q(k3[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[60]),
        .Q(k3[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[61]),
        .Q(k3[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[62]),
        .Q(k3[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[63]),
        .Q(k3[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[64] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[64]),
        .Q(k3[64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[65] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[65]),
        .Q(k3[65]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[66] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[66]),
        .Q(k3[66]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[67] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[67]),
        .Q(k3[67]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[68] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[68]),
        .Q(k3[68]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[69] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[69]),
        .Q(k3[69]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[6]),
        .Q(k3[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[70] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[70]),
        .Q(k3[70]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[71] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[71]),
        .Q(k3[71]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[72] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[72]),
        .Q(k3[72]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[73] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[73]),
        .Q(k3[73]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[74] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[74]),
        .Q(k3[74]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[75] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[75]),
        .Q(k3[75]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[76] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[76]),
        .Q(k3[76]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[77] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[77]),
        .Q(k3[77]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[78] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[78]),
        .Q(k3[78]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[79] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[79]),
        .Q(k3[79]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[7]),
        .Q(k3[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[80] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[80]),
        .Q(k3[80]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[81] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[81]),
        .Q(k3[81]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[82] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[82]),
        .Q(k3[82]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[83] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[83]),
        .Q(k3[83]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[84] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[84]),
        .Q(k3[84]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[85] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[85]),
        .Q(k3[85]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[86] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[86]),
        .Q(k3[86]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[87] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[87]),
        .Q(k3[87]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[88] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[88]),
        .Q(k3[88]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[89] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[89]),
        .Q(k3[89]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[8]),
        .Q(k3[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[90] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[90]),
        .Q(k3[90]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[91] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[91]),
        .Q(k3[91]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[92] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[92]),
        .Q(k3[92]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[93] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[93]),
        .Q(k3[93]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[94] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[94]),
        .Q(k3[94]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[95] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[95]),
        .Q(k3[95]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[96] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[96]),
        .Q(k3[96]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[97] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[97]),
        .Q(k3[97]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[98] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[98]),
        .Q(k3[98]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[99] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[99]),
        .Q(k3[99]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a3/out_1_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k2b[9]),
        .Q(k3[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_0/S_1/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \a4/S4_0/S_1/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,k3[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,k3[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\a4/S4_0/S_1/out_reg_n_0 ,\a4/S4_0/S_1/out_reg_n_1 ,\a4/S4_0/S_1/out_reg_n_2 ,\a4/S4_0/S_1/out_reg_n_3 ,\a4/S4_0/S_1/out_reg_n_4 ,\a4/S4_0/S_1/out_reg_n_5 ,\a4/S4_0/S_1/out_reg_n_6 ,\a4/S4_0/S_1/out_reg_n_7 ,\a4/k4a [23:16]}),
        .DOBDO({\a4/S4_0/S_1/out_reg_n_16 ,\a4/S4_0/S_1/out_reg_n_17 ,\a4/S4_0/S_1/out_reg_n_18 ,\a4/S4_0/S_1/out_reg_n_19 ,\a4/S4_0/S_1/out_reg_n_20 ,\a4/S4_0/S_1/out_reg_n_21 ,\a4/S4_0/S_1/out_reg_n_22 ,\a4/S4_0/S_1/out_reg_n_23 ,\a4/k4a [31:24]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_0/S_3/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \a4/S4_0/S_3/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,k3[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,k3[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\a4/S4_0/S_3/out_reg_n_0 ,\a4/S4_0/S_3/out_reg_n_1 ,\a4/S4_0/S_3/out_reg_n_2 ,\a4/S4_0/S_3/out_reg_n_3 ,\a4/S4_0/S_3/out_reg_n_4 ,\a4/S4_0/S_3/out_reg_n_5 ,\a4/S4_0/S_3/out_reg_n_6 ,\a4/S4_0/S_3/out_reg_n_7 ,\a4/k4a [7:0]}),
        .DOBDO({\a4/S4_0/S_3/out_reg_n_16 ,\a4/S4_0/S_3/out_reg_n_17 ,\a4/S4_0/S_3/out_reg_n_18 ,\a4/S4_0/S_3/out_reg_n_19 ,\a4/S4_0/S_3/out_reg_n_20 ,\a4/S4_0/S_3/out_reg_n_21 ,\a4/S4_0/S_3/out_reg_n_22 ,\a4/S4_0/S_3/out_reg_n_23 ,\a4/k4a [15:8]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[96]),
        .Q(\a4/k0a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[106]),
        .Q(\a4/k0a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[107]),
        .Q(\a4/k0a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[108]),
        .Q(\a4/k0a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[109]),
        .Q(\a4/k0a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[110]),
        .Q(\a4/k0a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[111]),
        .Q(\a4/k0a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[112]),
        .Q(\a4/k0a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[113]),
        .Q(\a4/k0a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[114]),
        .Q(\a4/k0a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[115]),
        .Q(\a4/k0a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[97]),
        .Q(\a4/k0a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[116]),
        .Q(\a4/k0a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[117]),
        .Q(\a4/k0a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[118]),
        .Q(\a4/k0a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[119]),
        .Q(\a4/k0a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[120]),
        .Q(\a4/k0a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[121]),
        .Q(\a4/k0a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[122]),
        .Q(\a4/k0a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v0 ),
        .Q(\a4/k0a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[124]),
        .Q(\a4/k0a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[125]),
        .Q(\a4/k0a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[98]),
        .Q(\a4/k0a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[126]),
        .Q(\a4/k0a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[127]),
        .Q(\a4/k0a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[99]),
        .Q(\a4/k0a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[100]),
        .Q(\a4/k0a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[101]),
        .Q(\a4/k0a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[102]),
        .Q(\a4/k0a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[103]),
        .Q(\a4/k0a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[104]),
        .Q(\a4/k0a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k0a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3[105]),
        .Q(\a4/k0a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [0]),
        .Q(\a4/k1a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [10]),
        .Q(\a4/k1a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [11]),
        .Q(\a4/k1a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [12]),
        .Q(\a4/k1a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [13]),
        .Q(\a4/k1a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [14]),
        .Q(\a4/k1a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [15]),
        .Q(\a4/k1a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [16]),
        .Q(\a4/k1a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [17]),
        .Q(\a4/k1a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [18]),
        .Q(\a4/k1a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [19]),
        .Q(\a4/k1a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [1]),
        .Q(\a4/k1a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [20]),
        .Q(\a4/k1a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [21]),
        .Q(\a4/k1a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [22]),
        .Q(\a4/k1a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [23]),
        .Q(\a4/k1a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [24]),
        .Q(\a4/k1a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [25]),
        .Q(\a4/k1a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [26]),
        .Q(\a4/k1a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\k1a[27]_i_1__2_n_0 ),
        .Q(\a4/k1a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [28]),
        .Q(\a4/k1a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [29]),
        .Q(\a4/k1a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [2]),
        .Q(\a4/k1a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [30]),
        .Q(\a4/k1a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [31]),
        .Q(\a4/k1a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [3]),
        .Q(\a4/k1a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [4]),
        .Q(\a4/k1a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [5]),
        .Q(\a4/k1a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [6]),
        .Q(\a4/k1a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [7]),
        .Q(\a4/k1a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [8]),
        .Q(\a4/k1a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k1a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v1 [9]),
        .Q(\a4/k1a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [0]),
        .Q(\a4/k2a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [10]),
        .Q(\a4/k2a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [11]),
        .Q(\a4/k2a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [12]),
        .Q(\a4/k2a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [13]),
        .Q(\a4/k2a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [14]),
        .Q(\a4/k2a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [15]),
        .Q(\a4/k2a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [16]),
        .Q(\a4/k2a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [17]),
        .Q(\a4/k2a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [18]),
        .Q(\a4/k2a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [19]),
        .Q(\a4/k2a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [1]),
        .Q(\a4/k2a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [20]),
        .Q(\a4/k2a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [21]),
        .Q(\a4/k2a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [22]),
        .Q(\a4/k2a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [23]),
        .Q(\a4/k2a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [24]),
        .Q(\a4/k2a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [25]),
        .Q(\a4/k2a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [26]),
        .Q(\a4/k2a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [27]),
        .Q(\a4/k2a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [28]),
        .Q(\a4/k2a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [29]),
        .Q(\a4/k2a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [2]),
        .Q(\a4/k2a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [30]),
        .Q(\a4/k2a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [31]),
        .Q(\a4/k2a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [3]),
        .Q(\a4/k2a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [4]),
        .Q(\a4/k2a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [5]),
        .Q(\a4/k2a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [6]),
        .Q(\a4/k2a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [7]),
        .Q(\a4/k2a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [8]),
        .Q(\a4/k2a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k2a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v2 [9]),
        .Q(\a4/k2a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [0]),
        .Q(\a4/k3a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [10]),
        .Q(\a4/k3a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [11]),
        .Q(\a4/k3a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [12]),
        .Q(\a4/k3a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [13]),
        .Q(\a4/k3a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [14]),
        .Q(\a4/k3a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [15]),
        .Q(\a4/k3a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [16]),
        .Q(\a4/k3a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [17]),
        .Q(\a4/k3a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [18]),
        .Q(\a4/k3a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [19]),
        .Q(\a4/k3a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [1]),
        .Q(\a4/k3a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [20]),
        .Q(\a4/k3a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [21]),
        .Q(\a4/k3a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [22]),
        .Q(\a4/k3a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [23]),
        .Q(\a4/k3a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [24]),
        .Q(\a4/k3a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [25]),
        .Q(\a4/k3a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [26]),
        .Q(\a4/k3a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [27]),
        .Q(\a4/k3a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [28]),
        .Q(\a4/k3a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [29]),
        .Q(\a4/k3a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [2]),
        .Q(\a4/k3a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [30]),
        .Q(\a4/k3a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [31]),
        .Q(\a4/k3a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [3]),
        .Q(\a4/k3a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [4]),
        .Q(\a4/k3a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [5]),
        .Q(\a4/k3a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [6]),
        .Q(\a4/k3a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [7]),
        .Q(\a4/k3a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [8]),
        .Q(\a4/k3a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/k3a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a4/v3 [9]),
        .Q(\a4/k3a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[0]),
        .Q(k4[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[100] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[100]),
        .Q(k4[100]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[101] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[101]),
        .Q(k4[101]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[102] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[102]),
        .Q(k4[102]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[103] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[103]),
        .Q(k4[103]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[104] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[104]),
        .Q(k4[104]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[105] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[105]),
        .Q(k4[105]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[106] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[106]),
        .Q(k4[106]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[107] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[107]),
        .Q(k4[107]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[108] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[108]),
        .Q(k4[108]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[109] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[109]),
        .Q(k4[109]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[10]),
        .Q(k4[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[110] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[110]),
        .Q(k4[110]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[111] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[111]),
        .Q(k4[111]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[112] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[112]),
        .Q(k4[112]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[113] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[113]),
        .Q(k4[113]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[114] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[114]),
        .Q(k4[114]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[115] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[115]),
        .Q(k4[115]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[116] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[116]),
        .Q(k4[116]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[117] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[117]),
        .Q(k4[117]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[118] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[118]),
        .Q(k4[118]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[119] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[119]),
        .Q(k4[119]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[11]),
        .Q(k4[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[120] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[120]),
        .Q(k4[120]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[121] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[121]),
        .Q(k4[121]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[122] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[122]),
        .Q(k4[122]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[123] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[123]),
        .Q(k4[123]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[124] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[124]),
        .Q(k4[124]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[125] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[125]),
        .Q(k4[125]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[126] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[126]),
        .Q(k4[126]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[127] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[127]),
        .Q(k4[127]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[12]),
        .Q(k4[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[13]),
        .Q(k4[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[14]),
        .Q(k4[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[15]),
        .Q(k4[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[16]),
        .Q(k4[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[17]),
        .Q(k4[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[18]),
        .Q(k4[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[19]),
        .Q(k4[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[1]),
        .Q(k4[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[20]),
        .Q(k4[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[21]),
        .Q(k4[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[22]),
        .Q(k4[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[23]),
        .Q(k4[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[24]),
        .Q(k4[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[25]),
        .Q(k4[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[26]),
        .Q(k4[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[27]),
        .Q(k4[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[28]),
        .Q(k4[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[29]),
        .Q(k4[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[2]),
        .Q(k4[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[30]),
        .Q(k4[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[31]),
        .Q(k4[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[32]),
        .Q(k4[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[33]),
        .Q(k4[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[34]),
        .Q(k4[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[35]),
        .Q(k4[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[36]),
        .Q(k4[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[37]),
        .Q(k4[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[38]),
        .Q(k4[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[39]),
        .Q(k4[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[3]),
        .Q(k4[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[40]),
        .Q(k4[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[41]),
        .Q(k4[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[42]),
        .Q(k4[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[43]),
        .Q(k4[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[44]),
        .Q(k4[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[45]),
        .Q(k4[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[46]),
        .Q(k4[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[47]),
        .Q(k4[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[48]),
        .Q(k4[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[49]),
        .Q(k4[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[4]),
        .Q(k4[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[50]),
        .Q(k4[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[51]),
        .Q(k4[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[52]),
        .Q(k4[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[53]),
        .Q(k4[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[54]),
        .Q(k4[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[55]),
        .Q(k4[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[56]),
        .Q(k4[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[57]),
        .Q(k4[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[58]),
        .Q(k4[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[59]),
        .Q(k4[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[5]),
        .Q(k4[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[60]),
        .Q(k4[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[61]),
        .Q(k4[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[62]),
        .Q(k4[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[63]),
        .Q(k4[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[64] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[64]),
        .Q(k4[64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[65] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[65]),
        .Q(k4[65]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[66] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[66]),
        .Q(k4[66]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[67] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[67]),
        .Q(k4[67]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[68] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[68]),
        .Q(k4[68]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[69] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[69]),
        .Q(k4[69]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[6]),
        .Q(k4[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[70] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[70]),
        .Q(k4[70]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[71] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[71]),
        .Q(k4[71]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[72] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[72]),
        .Q(k4[72]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[73] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[73]),
        .Q(k4[73]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[74] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[74]),
        .Q(k4[74]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[75] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[75]),
        .Q(k4[75]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[76] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[76]),
        .Q(k4[76]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[77] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[77]),
        .Q(k4[77]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[78] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[78]),
        .Q(k4[78]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[79] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[79]),
        .Q(k4[79]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[7]),
        .Q(k4[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[80] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[80]),
        .Q(k4[80]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[81] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[81]),
        .Q(k4[81]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[82] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[82]),
        .Q(k4[82]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[83] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[83]),
        .Q(k4[83]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[84] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[84]),
        .Q(k4[84]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[85] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[85]),
        .Q(k4[85]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[86] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[86]),
        .Q(k4[86]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[87] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[87]),
        .Q(k4[87]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[88] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[88]),
        .Q(k4[88]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[89] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[89]),
        .Q(k4[89]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[8]),
        .Q(k4[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[90] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[90]),
        .Q(k4[90]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[91] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[91]),
        .Q(k4[91]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[92] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[92]),
        .Q(k4[92]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[93] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[93]),
        .Q(k4[93]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[94] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[94]),
        .Q(k4[94]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[95] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[95]),
        .Q(k4[95]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[96] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[96]),
        .Q(k4[96]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[97] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[97]),
        .Q(k4[97]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[98] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[98]),
        .Q(k4[98]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[99] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[99]),
        .Q(k4[99]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a4/out_1_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k3b[9]),
        .Q(k4[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_0/S_1/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \a5/S4_0/S_1/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,k4[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,k4[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\a5/S4_0/S_1/out_reg_n_0 ,\a5/S4_0/S_1/out_reg_n_1 ,\a5/S4_0/S_1/out_reg_n_2 ,\a5/S4_0/S_1/out_reg_n_3 ,\a5/S4_0/S_1/out_reg_n_4 ,\a5/S4_0/S_1/out_reg_n_5 ,\a5/S4_0/S_1/out_reg_n_6 ,\a5/S4_0/S_1/out_reg_n_7 ,\a5/k4a [23:16]}),
        .DOBDO({\a5/S4_0/S_1/out_reg_n_16 ,\a5/S4_0/S_1/out_reg_n_17 ,\a5/S4_0/S_1/out_reg_n_18 ,\a5/S4_0/S_1/out_reg_n_19 ,\a5/S4_0/S_1/out_reg_n_20 ,\a5/S4_0/S_1/out_reg_n_21 ,\a5/S4_0/S_1/out_reg_n_22 ,\a5/S4_0/S_1/out_reg_n_23 ,\a5/k4a [31:24]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_0/S_3/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \a5/S4_0/S_3/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,k4[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,k4[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\a5/S4_0/S_3/out_reg_n_0 ,\a5/S4_0/S_3/out_reg_n_1 ,\a5/S4_0/S_3/out_reg_n_2 ,\a5/S4_0/S_3/out_reg_n_3 ,\a5/S4_0/S_3/out_reg_n_4 ,\a5/S4_0/S_3/out_reg_n_5 ,\a5/S4_0/S_3/out_reg_n_6 ,\a5/S4_0/S_3/out_reg_n_7 ,\a5/k4a [7:0]}),
        .DOBDO({\a5/S4_0/S_3/out_reg_n_16 ,\a5/S4_0/S_3/out_reg_n_17 ,\a5/S4_0/S_3/out_reg_n_18 ,\a5/S4_0/S_3/out_reg_n_19 ,\a5/S4_0/S_3/out_reg_n_20 ,\a5/S4_0/S_3/out_reg_n_21 ,\a5/S4_0/S_3/out_reg_n_22 ,\a5/S4_0/S_3/out_reg_n_23 ,\a5/k4a [15:8]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[96]),
        .Q(\a5/k0a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[106]),
        .Q(\a5/k0a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[107]),
        .Q(\a5/k0a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[108]),
        .Q(\a5/k0a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[109]),
        .Q(\a5/k0a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[110]),
        .Q(\a5/k0a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[111]),
        .Q(\a5/k0a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[112]),
        .Q(\a5/k0a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[113]),
        .Q(\a5/k0a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[114]),
        .Q(\a5/k0a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[115]),
        .Q(\a5/k0a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[97]),
        .Q(\a5/k0a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[116]),
        .Q(\a5/k0a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[117]),
        .Q(\a5/k0a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[118]),
        .Q(\a5/k0a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[119]),
        .Q(\a5/k0a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[120]),
        .Q(\a5/k0a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[121]),
        .Q(\a5/k0a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[122]),
        .Q(\a5/k0a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[123]),
        .Q(\a5/k0a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v0 ),
        .Q(\a5/k0a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[125]),
        .Q(\a5/k0a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[98]),
        .Q(\a5/k0a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[126]),
        .Q(\a5/k0a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[127]),
        .Q(\a5/k0a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[99]),
        .Q(\a5/k0a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[100]),
        .Q(\a5/k0a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[101]),
        .Q(\a5/k0a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[102]),
        .Q(\a5/k0a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[103]),
        .Q(\a5/k0a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[104]),
        .Q(\a5/k0a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k0a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4[105]),
        .Q(\a5/k0a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [0]),
        .Q(\a5/k1a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [10]),
        .Q(\a5/k1a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [11]),
        .Q(\a5/k1a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [12]),
        .Q(\a5/k1a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [13]),
        .Q(\a5/k1a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [14]),
        .Q(\a5/k1a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [15]),
        .Q(\a5/k1a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [16]),
        .Q(\a5/k1a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [17]),
        .Q(\a5/k1a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [18]),
        .Q(\a5/k1a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [19]),
        .Q(\a5/k1a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [1]),
        .Q(\a5/k1a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [20]),
        .Q(\a5/k1a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [21]),
        .Q(\a5/k1a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [22]),
        .Q(\a5/k1a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [23]),
        .Q(\a5/k1a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [24]),
        .Q(\a5/k1a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [25]),
        .Q(\a5/k1a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [26]),
        .Q(\a5/k1a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [27]),
        .Q(\a5/k1a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\k1a[28]_i_1__3_n_0 ),
        .Q(\a5/k1a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [29]),
        .Q(\a5/k1a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [2]),
        .Q(\a5/k1a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [30]),
        .Q(\a5/k1a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [31]),
        .Q(\a5/k1a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [3]),
        .Q(\a5/k1a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [4]),
        .Q(\a5/k1a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [5]),
        .Q(\a5/k1a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [6]),
        .Q(\a5/k1a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [7]),
        .Q(\a5/k1a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [8]),
        .Q(\a5/k1a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k1a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v1 [9]),
        .Q(\a5/k1a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [0]),
        .Q(\a5/k2a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [10]),
        .Q(\a5/k2a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [11]),
        .Q(\a5/k2a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [12]),
        .Q(\a5/k2a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [13]),
        .Q(\a5/k2a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [14]),
        .Q(\a5/k2a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [15]),
        .Q(\a5/k2a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [16]),
        .Q(\a5/k2a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [17]),
        .Q(\a5/k2a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [18]),
        .Q(\a5/k2a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [19]),
        .Q(\a5/k2a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [1]),
        .Q(\a5/k2a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [20]),
        .Q(\a5/k2a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [21]),
        .Q(\a5/k2a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [22]),
        .Q(\a5/k2a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [23]),
        .Q(\a5/k2a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [24]),
        .Q(\a5/k2a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [25]),
        .Q(\a5/k2a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [26]),
        .Q(\a5/k2a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [27]),
        .Q(\a5/k2a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [28]),
        .Q(\a5/k2a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [29]),
        .Q(\a5/k2a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [2]),
        .Q(\a5/k2a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [30]),
        .Q(\a5/k2a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [31]),
        .Q(\a5/k2a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [3]),
        .Q(\a5/k2a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [4]),
        .Q(\a5/k2a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [5]),
        .Q(\a5/k2a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [6]),
        .Q(\a5/k2a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [7]),
        .Q(\a5/k2a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [8]),
        .Q(\a5/k2a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k2a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v2 [9]),
        .Q(\a5/k2a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [0]),
        .Q(\a5/k3a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [10]),
        .Q(\a5/k3a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [11]),
        .Q(\a5/k3a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [12]),
        .Q(\a5/k3a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [13]),
        .Q(\a5/k3a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [14]),
        .Q(\a5/k3a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [15]),
        .Q(\a5/k3a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [16]),
        .Q(\a5/k3a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [17]),
        .Q(\a5/k3a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [18]),
        .Q(\a5/k3a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [19]),
        .Q(\a5/k3a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [1]),
        .Q(\a5/k3a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [20]),
        .Q(\a5/k3a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [21]),
        .Q(\a5/k3a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [22]),
        .Q(\a5/k3a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [23]),
        .Q(\a5/k3a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [24]),
        .Q(\a5/k3a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [25]),
        .Q(\a5/k3a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [26]),
        .Q(\a5/k3a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [27]),
        .Q(\a5/k3a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [28]),
        .Q(\a5/k3a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [29]),
        .Q(\a5/k3a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [2]),
        .Q(\a5/k3a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [30]),
        .Q(\a5/k3a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [31]),
        .Q(\a5/k3a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [3]),
        .Q(\a5/k3a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [4]),
        .Q(\a5/k3a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [5]),
        .Q(\a5/k3a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [6]),
        .Q(\a5/k3a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [7]),
        .Q(\a5/k3a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [8]),
        .Q(\a5/k3a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/k3a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a5/v3 [9]),
        .Q(\a5/k3a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[0]),
        .Q(k5[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[100] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[100]),
        .Q(k5[100]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[101] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[101]),
        .Q(k5[101]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[102] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[102]),
        .Q(k5[102]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[103] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[103]),
        .Q(k5[103]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[104] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[104]),
        .Q(k5[104]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[105] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[105]),
        .Q(k5[105]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[106] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[106]),
        .Q(k5[106]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[107] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[107]),
        .Q(k5[107]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[108] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[108]),
        .Q(k5[108]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[109] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[109]),
        .Q(k5[109]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[10]),
        .Q(k5[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[110] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[110]),
        .Q(k5[110]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[111] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[111]),
        .Q(k5[111]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[112] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[112]),
        .Q(k5[112]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[113] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[113]),
        .Q(k5[113]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[114] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[114]),
        .Q(k5[114]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[115] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[115]),
        .Q(k5[115]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[116] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[116]),
        .Q(k5[116]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[117] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[117]),
        .Q(k5[117]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[118] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[118]),
        .Q(k5[118]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[119] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[119]),
        .Q(k5[119]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[11]),
        .Q(k5[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[120] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[120]),
        .Q(k5[120]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[121] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[121]),
        .Q(k5[121]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[122] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[122]),
        .Q(k5[122]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[123] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[123]),
        .Q(k5[123]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[124] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[124]),
        .Q(k5[124]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[125] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[125]),
        .Q(k5[125]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[126] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[126]),
        .Q(k5[126]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[127] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[127]),
        .Q(k5[127]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[12]),
        .Q(k5[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[13]),
        .Q(k5[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[14]),
        .Q(k5[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[15]),
        .Q(k5[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[16]),
        .Q(k5[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[17]),
        .Q(k5[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[18]),
        .Q(k5[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[19]),
        .Q(k5[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[1]),
        .Q(k5[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[20]),
        .Q(k5[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[21]),
        .Q(k5[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[22]),
        .Q(k5[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[23]),
        .Q(k5[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[24]),
        .Q(k5[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[25]),
        .Q(k5[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[26]),
        .Q(k5[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[27]),
        .Q(k5[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[28]),
        .Q(k5[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[29]),
        .Q(k5[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[2]),
        .Q(k5[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[30]),
        .Q(k5[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[31]),
        .Q(k5[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[32]),
        .Q(k5[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[33]),
        .Q(k5[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[34]),
        .Q(k5[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[35]),
        .Q(k5[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[36]),
        .Q(k5[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[37]),
        .Q(k5[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[38]),
        .Q(k5[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[39]),
        .Q(k5[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[3]),
        .Q(k5[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[40]),
        .Q(k5[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[41]),
        .Q(k5[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[42]),
        .Q(k5[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[43]),
        .Q(k5[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[44]),
        .Q(k5[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[45]),
        .Q(k5[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[46]),
        .Q(k5[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[47]),
        .Q(k5[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[48]),
        .Q(k5[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[49]),
        .Q(k5[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[4]),
        .Q(k5[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[50]),
        .Q(k5[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[51]),
        .Q(k5[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[52]),
        .Q(k5[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[53]),
        .Q(k5[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[54]),
        .Q(k5[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[55]),
        .Q(k5[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[56]),
        .Q(k5[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[57]),
        .Q(k5[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[58]),
        .Q(k5[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[59]),
        .Q(k5[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[5]),
        .Q(k5[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[60]),
        .Q(k5[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[61]),
        .Q(k5[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[62]),
        .Q(k5[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[63]),
        .Q(k5[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[64] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[64]),
        .Q(k5[64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[65] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[65]),
        .Q(k5[65]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[66] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[66]),
        .Q(k5[66]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[67] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[67]),
        .Q(k5[67]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[68] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[68]),
        .Q(k5[68]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[69] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[69]),
        .Q(k5[69]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[6]),
        .Q(k5[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[70] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[70]),
        .Q(k5[70]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[71] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[71]),
        .Q(k5[71]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[72] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[72]),
        .Q(k5[72]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[73] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[73]),
        .Q(k5[73]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[74] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[74]),
        .Q(k5[74]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[75] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[75]),
        .Q(k5[75]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[76] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[76]),
        .Q(k5[76]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[77] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[77]),
        .Q(k5[77]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[78] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[78]),
        .Q(k5[78]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[79] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[79]),
        .Q(k5[79]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[7]),
        .Q(k5[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[80] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[80]),
        .Q(k5[80]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[81] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[81]),
        .Q(k5[81]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[82] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[82]),
        .Q(k5[82]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[83] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[83]),
        .Q(k5[83]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[84] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[84]),
        .Q(k5[84]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[85] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[85]),
        .Q(k5[85]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[86] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[86]),
        .Q(k5[86]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[87] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[87]),
        .Q(k5[87]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[88] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[88]),
        .Q(k5[88]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[89] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[89]),
        .Q(k5[89]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[8]),
        .Q(k5[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[90] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[90]),
        .Q(k5[90]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[91] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[91]),
        .Q(k5[91]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[92] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[92]),
        .Q(k5[92]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[93] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[93]),
        .Q(k5[93]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[94] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[94]),
        .Q(k5[94]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[95] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[95]),
        .Q(k5[95]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[96] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[96]),
        .Q(k5[96]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[97] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[97]),
        .Q(k5[97]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[98] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[98]),
        .Q(k5[98]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[99] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[99]),
        .Q(k5[99]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a5/out_1_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k4b[9]),
        .Q(k5[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_0/S_1/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \a6/S4_0/S_1/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,k5[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,k5[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\a6/S4_0/S_1/out_reg_n_0 ,\a6/S4_0/S_1/out_reg_n_1 ,\a6/S4_0/S_1/out_reg_n_2 ,\a6/S4_0/S_1/out_reg_n_3 ,\a6/S4_0/S_1/out_reg_n_4 ,\a6/S4_0/S_1/out_reg_n_5 ,\a6/S4_0/S_1/out_reg_n_6 ,\a6/S4_0/S_1/out_reg_n_7 ,\a6/k4a [23:16]}),
        .DOBDO({\a6/S4_0/S_1/out_reg_n_16 ,\a6/S4_0/S_1/out_reg_n_17 ,\a6/S4_0/S_1/out_reg_n_18 ,\a6/S4_0/S_1/out_reg_n_19 ,\a6/S4_0/S_1/out_reg_n_20 ,\a6/S4_0/S_1/out_reg_n_21 ,\a6/S4_0/S_1/out_reg_n_22 ,\a6/S4_0/S_1/out_reg_n_23 ,\a6/k4a [31:24]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_0/S_3/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \a6/S4_0/S_3/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,k5[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,k5[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\a6/S4_0/S_3/out_reg_n_0 ,\a6/S4_0/S_3/out_reg_n_1 ,\a6/S4_0/S_3/out_reg_n_2 ,\a6/S4_0/S_3/out_reg_n_3 ,\a6/S4_0/S_3/out_reg_n_4 ,\a6/S4_0/S_3/out_reg_n_5 ,\a6/S4_0/S_3/out_reg_n_6 ,\a6/S4_0/S_3/out_reg_n_7 ,\a6/k4a [7:0]}),
        .DOBDO({\a6/S4_0/S_3/out_reg_n_16 ,\a6/S4_0/S_3/out_reg_n_17 ,\a6/S4_0/S_3/out_reg_n_18 ,\a6/S4_0/S_3/out_reg_n_19 ,\a6/S4_0/S_3/out_reg_n_20 ,\a6/S4_0/S_3/out_reg_n_21 ,\a6/S4_0/S_3/out_reg_n_22 ,\a6/S4_0/S_3/out_reg_n_23 ,\a6/k4a [15:8]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[96]),
        .Q(\a6/k0a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[106]),
        .Q(\a6/k0a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[107]),
        .Q(\a6/k0a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[108]),
        .Q(\a6/k0a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[109]),
        .Q(\a6/k0a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[110]),
        .Q(\a6/k0a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[111]),
        .Q(\a6/k0a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[112]),
        .Q(\a6/k0a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[113]),
        .Q(\a6/k0a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[114]),
        .Q(\a6/k0a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[115]),
        .Q(\a6/k0a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[97]),
        .Q(\a6/k0a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[116]),
        .Q(\a6/k0a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[117]),
        .Q(\a6/k0a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[118]),
        .Q(\a6/k0a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[119]),
        .Q(\a6/k0a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[120]),
        .Q(\a6/k0a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[121]),
        .Q(\a6/k0a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[122]),
        .Q(\a6/k0a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[123]),
        .Q(\a6/k0a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[124]),
        .Q(\a6/k0a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v0 ),
        .Q(\a6/k0a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[98]),
        .Q(\a6/k0a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[126]),
        .Q(\a6/k0a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[127]),
        .Q(\a6/k0a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[99]),
        .Q(\a6/k0a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[100]),
        .Q(\a6/k0a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[101]),
        .Q(\a6/k0a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[102]),
        .Q(\a6/k0a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[103]),
        .Q(\a6/k0a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[104]),
        .Q(\a6/k0a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k0a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5[105]),
        .Q(\a6/k0a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [0]),
        .Q(\a6/k1a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [10]),
        .Q(\a6/k1a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [11]),
        .Q(\a6/k1a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [12]),
        .Q(\a6/k1a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [13]),
        .Q(\a6/k1a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [14]),
        .Q(\a6/k1a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [15]),
        .Q(\a6/k1a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [16]),
        .Q(\a6/k1a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [17]),
        .Q(\a6/k1a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [18]),
        .Q(\a6/k1a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [19]),
        .Q(\a6/k1a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [1]),
        .Q(\a6/k1a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [20]),
        .Q(\a6/k1a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [21]),
        .Q(\a6/k1a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [22]),
        .Q(\a6/k1a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [23]),
        .Q(\a6/k1a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [24]),
        .Q(\a6/k1a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [25]),
        .Q(\a6/k1a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [26]),
        .Q(\a6/k1a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [27]),
        .Q(\a6/k1a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [28]),
        .Q(\a6/k1a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\k1a[29]_i_1__4_n_0 ),
        .Q(\a6/k1a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [2]),
        .Q(\a6/k1a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [30]),
        .Q(\a6/k1a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [31]),
        .Q(\a6/k1a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [3]),
        .Q(\a6/k1a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [4]),
        .Q(\a6/k1a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [5]),
        .Q(\a6/k1a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [6]),
        .Q(\a6/k1a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [7]),
        .Q(\a6/k1a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [8]),
        .Q(\a6/k1a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k1a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v1 [9]),
        .Q(\a6/k1a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [0]),
        .Q(\a6/k2a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [10]),
        .Q(\a6/k2a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [11]),
        .Q(\a6/k2a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [12]),
        .Q(\a6/k2a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [13]),
        .Q(\a6/k2a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [14]),
        .Q(\a6/k2a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [15]),
        .Q(\a6/k2a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [16]),
        .Q(\a6/k2a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [17]),
        .Q(\a6/k2a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [18]),
        .Q(\a6/k2a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [19]),
        .Q(\a6/k2a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [1]),
        .Q(\a6/k2a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [20]),
        .Q(\a6/k2a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [21]),
        .Q(\a6/k2a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [22]),
        .Q(\a6/k2a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [23]),
        .Q(\a6/k2a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [24]),
        .Q(\a6/k2a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [25]),
        .Q(\a6/k2a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [26]),
        .Q(\a6/k2a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [27]),
        .Q(\a6/k2a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [28]),
        .Q(\a6/k2a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [29]),
        .Q(\a6/k2a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [2]),
        .Q(\a6/k2a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [30]),
        .Q(\a6/k2a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [31]),
        .Q(\a6/k2a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [3]),
        .Q(\a6/k2a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [4]),
        .Q(\a6/k2a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [5]),
        .Q(\a6/k2a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [6]),
        .Q(\a6/k2a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [7]),
        .Q(\a6/k2a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [8]),
        .Q(\a6/k2a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k2a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v2 [9]),
        .Q(\a6/k2a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [0]),
        .Q(\a6/k3a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [10]),
        .Q(\a6/k3a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [11]),
        .Q(\a6/k3a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [12]),
        .Q(\a6/k3a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [13]),
        .Q(\a6/k3a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [14]),
        .Q(\a6/k3a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [15]),
        .Q(\a6/k3a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [16]),
        .Q(\a6/k3a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [17]),
        .Q(\a6/k3a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [18]),
        .Q(\a6/k3a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [19]),
        .Q(\a6/k3a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [1]),
        .Q(\a6/k3a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [20]),
        .Q(\a6/k3a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [21]),
        .Q(\a6/k3a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [22]),
        .Q(\a6/k3a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [23]),
        .Q(\a6/k3a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [24]),
        .Q(\a6/k3a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [25]),
        .Q(\a6/k3a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [26]),
        .Q(\a6/k3a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [27]),
        .Q(\a6/k3a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [28]),
        .Q(\a6/k3a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [29]),
        .Q(\a6/k3a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [2]),
        .Q(\a6/k3a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [30]),
        .Q(\a6/k3a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [31]),
        .Q(\a6/k3a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [3]),
        .Q(\a6/k3a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [4]),
        .Q(\a6/k3a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [5]),
        .Q(\a6/k3a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [6]),
        .Q(\a6/k3a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [7]),
        .Q(\a6/k3a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [8]),
        .Q(\a6/k3a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/k3a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a6/v3 [9]),
        .Q(\a6/k3a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[0]),
        .Q(k6[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[100] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[100]),
        .Q(k6[100]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[101] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[101]),
        .Q(k6[101]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[102] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[102]),
        .Q(k6[102]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[103] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[103]),
        .Q(k6[103]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[104] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[104]),
        .Q(k6[104]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[105] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[105]),
        .Q(k6[105]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[106] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[106]),
        .Q(k6[106]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[107] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[107]),
        .Q(k6[107]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[108] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[108]),
        .Q(k6[108]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[109] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[109]),
        .Q(k6[109]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[10]),
        .Q(k6[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[110] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[110]),
        .Q(k6[110]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[111] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[111]),
        .Q(k6[111]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[112] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[112]),
        .Q(k6[112]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[113] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[113]),
        .Q(k6[113]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[114] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[114]),
        .Q(k6[114]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[115] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[115]),
        .Q(k6[115]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[116] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[116]),
        .Q(k6[116]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[117] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[117]),
        .Q(k6[117]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[118] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[118]),
        .Q(k6[118]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[119] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[119]),
        .Q(k6[119]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[11]),
        .Q(k6[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[120] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[120]),
        .Q(k6[120]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[121] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[121]),
        .Q(k6[121]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[122] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[122]),
        .Q(k6[122]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[123] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[123]),
        .Q(k6[123]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[124] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[124]),
        .Q(k6[124]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[125] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[125]),
        .Q(k6[125]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[126] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[126]),
        .Q(k6[126]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[127] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[127]),
        .Q(k6[127]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[12]),
        .Q(k6[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[13]),
        .Q(k6[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[14]),
        .Q(k6[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[15]),
        .Q(k6[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[16]),
        .Q(k6[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[17]),
        .Q(k6[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[18]),
        .Q(k6[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[19]),
        .Q(k6[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[1]),
        .Q(k6[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[20]),
        .Q(k6[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[21]),
        .Q(k6[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[22]),
        .Q(k6[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[23]),
        .Q(k6[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[24]),
        .Q(k6[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[25]),
        .Q(k6[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[26]),
        .Q(k6[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[27]),
        .Q(k6[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[28]),
        .Q(k6[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[29]),
        .Q(k6[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[2]),
        .Q(k6[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[30]),
        .Q(k6[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[31]),
        .Q(k6[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[32]),
        .Q(k6[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[33]),
        .Q(k6[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[34]),
        .Q(k6[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[35]),
        .Q(k6[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[36]),
        .Q(k6[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[37]),
        .Q(k6[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[38]),
        .Q(k6[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[39]),
        .Q(k6[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[3]),
        .Q(k6[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[40]),
        .Q(k6[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[41]),
        .Q(k6[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[42]),
        .Q(k6[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[43]),
        .Q(k6[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[44]),
        .Q(k6[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[45]),
        .Q(k6[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[46]),
        .Q(k6[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[47]),
        .Q(k6[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[48]),
        .Q(k6[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[49]),
        .Q(k6[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[4]),
        .Q(k6[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[50]),
        .Q(k6[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[51]),
        .Q(k6[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[52]),
        .Q(k6[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[53]),
        .Q(k6[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[54]),
        .Q(k6[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[55]),
        .Q(k6[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[56]),
        .Q(k6[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[57]),
        .Q(k6[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[58]),
        .Q(k6[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[59]),
        .Q(k6[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[5]),
        .Q(k6[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[60]),
        .Q(k6[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[61]),
        .Q(k6[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[62]),
        .Q(k6[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[63]),
        .Q(k6[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[64] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[64]),
        .Q(k6[64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[65] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[65]),
        .Q(k6[65]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[66] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[66]),
        .Q(k6[66]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[67] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[67]),
        .Q(k6[67]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[68] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[68]),
        .Q(k6[68]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[69] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[69]),
        .Q(k6[69]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[6]),
        .Q(k6[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[70] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[70]),
        .Q(k6[70]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[71] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[71]),
        .Q(k6[71]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[72] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[72]),
        .Q(k6[72]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[73] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[73]),
        .Q(k6[73]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[74] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[74]),
        .Q(k6[74]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[75] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[75]),
        .Q(k6[75]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[76] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[76]),
        .Q(k6[76]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[77] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[77]),
        .Q(k6[77]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[78] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[78]),
        .Q(k6[78]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[79] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[79]),
        .Q(k6[79]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[7]),
        .Q(k6[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[80] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[80]),
        .Q(k6[80]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[81] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[81]),
        .Q(k6[81]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[82] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[82]),
        .Q(k6[82]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[83] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[83]),
        .Q(k6[83]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[84] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[84]),
        .Q(k6[84]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[85] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[85]),
        .Q(k6[85]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[86] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[86]),
        .Q(k6[86]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[87] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[87]),
        .Q(k6[87]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[88] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[88]),
        .Q(k6[88]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[89] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[89]),
        .Q(k6[89]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[8]),
        .Q(k6[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[90] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[90]),
        .Q(k6[90]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[91] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[91]),
        .Q(k6[91]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[92] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[92]),
        .Q(k6[92]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[93] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[93]),
        .Q(k6[93]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[94] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[94]),
        .Q(k6[94]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[95] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[95]),
        .Q(k6[95]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[96] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[96]),
        .Q(k6[96]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[97] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[97]),
        .Q(k6[97]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[98] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[98]),
        .Q(k6[98]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[99] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[99]),
        .Q(k6[99]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a6/out_1_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k5b[9]),
        .Q(k6[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_0/S_1/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \a7/S4_0/S_1/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,k6[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,k6[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\a7/S4_0/S_1/out_reg_n_0 ,\a7/S4_0/S_1/out_reg_n_1 ,\a7/S4_0/S_1/out_reg_n_2 ,\a7/S4_0/S_1/out_reg_n_3 ,\a7/S4_0/S_1/out_reg_n_4 ,\a7/S4_0/S_1/out_reg_n_5 ,\a7/S4_0/S_1/out_reg_n_6 ,\a7/S4_0/S_1/out_reg_n_7 ,\a7/k4a [23:16]}),
        .DOBDO({\a7/S4_0/S_1/out_reg_n_16 ,\a7/S4_0/S_1/out_reg_n_17 ,\a7/S4_0/S_1/out_reg_n_18 ,\a7/S4_0/S_1/out_reg_n_19 ,\a7/S4_0/S_1/out_reg_n_20 ,\a7/S4_0/S_1/out_reg_n_21 ,\a7/S4_0/S_1/out_reg_n_22 ,\a7/S4_0/S_1/out_reg_n_23 ,\a7/k4a [31:24]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_0/S_3/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \a7/S4_0/S_3/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,k6[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,k6[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\a7/S4_0/S_3/out_reg_n_0 ,\a7/S4_0/S_3/out_reg_n_1 ,\a7/S4_0/S_3/out_reg_n_2 ,\a7/S4_0/S_3/out_reg_n_3 ,\a7/S4_0/S_3/out_reg_n_4 ,\a7/S4_0/S_3/out_reg_n_5 ,\a7/S4_0/S_3/out_reg_n_6 ,\a7/S4_0/S_3/out_reg_n_7 ,\a7/k4a [7:0]}),
        .DOBDO({\a7/S4_0/S_3/out_reg_n_16 ,\a7/S4_0/S_3/out_reg_n_17 ,\a7/S4_0/S_3/out_reg_n_18 ,\a7/S4_0/S_3/out_reg_n_19 ,\a7/S4_0/S_3/out_reg_n_20 ,\a7/S4_0/S_3/out_reg_n_21 ,\a7/S4_0/S_3/out_reg_n_22 ,\a7/S4_0/S_3/out_reg_n_23 ,\a7/k4a [15:8]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[96]),
        .Q(\a7/k0a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[106]),
        .Q(\a7/k0a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[107]),
        .Q(\a7/k0a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[108]),
        .Q(\a7/k0a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[109]),
        .Q(\a7/k0a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[110]),
        .Q(\a7/k0a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[111]),
        .Q(\a7/k0a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[112]),
        .Q(\a7/k0a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[113]),
        .Q(\a7/k0a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[114]),
        .Q(\a7/k0a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[115]),
        .Q(\a7/k0a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[97]),
        .Q(\a7/k0a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[116]),
        .Q(\a7/k0a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[117]),
        .Q(\a7/k0a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[118]),
        .Q(\a7/k0a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[119]),
        .Q(\a7/k0a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[120]),
        .Q(\a7/k0a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[121]),
        .Q(\a7/k0a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[122]),
        .Q(\a7/k0a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[123]),
        .Q(\a7/k0a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[124]),
        .Q(\a7/k0a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[125]),
        .Q(\a7/k0a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[98]),
        .Q(\a7/k0a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v0 ),
        .Q(\a7/k0a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[127]),
        .Q(\a7/k0a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[99]),
        .Q(\a7/k0a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[100]),
        .Q(\a7/k0a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[101]),
        .Q(\a7/k0a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[102]),
        .Q(\a7/k0a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[103]),
        .Q(\a7/k0a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[104]),
        .Q(\a7/k0a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k0a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6[105]),
        .Q(\a7/k0a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [0]),
        .Q(\a7/k1a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [10]),
        .Q(\a7/k1a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [11]),
        .Q(\a7/k1a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [12]),
        .Q(\a7/k1a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [13]),
        .Q(\a7/k1a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [14]),
        .Q(\a7/k1a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [15]),
        .Q(\a7/k1a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [16]),
        .Q(\a7/k1a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [17]),
        .Q(\a7/k1a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [18]),
        .Q(\a7/k1a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [19]),
        .Q(\a7/k1a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [1]),
        .Q(\a7/k1a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [20]),
        .Q(\a7/k1a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [21]),
        .Q(\a7/k1a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [22]),
        .Q(\a7/k1a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [23]),
        .Q(\a7/k1a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [24]),
        .Q(\a7/k1a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [25]),
        .Q(\a7/k1a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [26]),
        .Q(\a7/k1a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [27]),
        .Q(\a7/k1a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [28]),
        .Q(\a7/k1a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [29]),
        .Q(\a7/k1a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [2]),
        .Q(\a7/k1a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\k1a[30]_i_1__5_n_0 ),
        .Q(\a7/k1a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [31]),
        .Q(\a7/k1a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [3]),
        .Q(\a7/k1a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [4]),
        .Q(\a7/k1a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [5]),
        .Q(\a7/k1a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [6]),
        .Q(\a7/k1a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [7]),
        .Q(\a7/k1a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [8]),
        .Q(\a7/k1a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k1a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v1 [9]),
        .Q(\a7/k1a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [0]),
        .Q(\a7/k2a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [10]),
        .Q(\a7/k2a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [11]),
        .Q(\a7/k2a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [12]),
        .Q(\a7/k2a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [13]),
        .Q(\a7/k2a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [14]),
        .Q(\a7/k2a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [15]),
        .Q(\a7/k2a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [16]),
        .Q(\a7/k2a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [17]),
        .Q(\a7/k2a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [18]),
        .Q(\a7/k2a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [19]),
        .Q(\a7/k2a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [1]),
        .Q(\a7/k2a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [20]),
        .Q(\a7/k2a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [21]),
        .Q(\a7/k2a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [22]),
        .Q(\a7/k2a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [23]),
        .Q(\a7/k2a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [24]),
        .Q(\a7/k2a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [25]),
        .Q(\a7/k2a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [26]),
        .Q(\a7/k2a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [27]),
        .Q(\a7/k2a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [28]),
        .Q(\a7/k2a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [29]),
        .Q(\a7/k2a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [2]),
        .Q(\a7/k2a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [30]),
        .Q(\a7/k2a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [31]),
        .Q(\a7/k2a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [3]),
        .Q(\a7/k2a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [4]),
        .Q(\a7/k2a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [5]),
        .Q(\a7/k2a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [6]),
        .Q(\a7/k2a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [7]),
        .Q(\a7/k2a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [8]),
        .Q(\a7/k2a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k2a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v2 [9]),
        .Q(\a7/k2a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [0]),
        .Q(\a7/k3a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [10]),
        .Q(\a7/k3a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [11]),
        .Q(\a7/k3a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [12]),
        .Q(\a7/k3a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [13]),
        .Q(\a7/k3a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [14]),
        .Q(\a7/k3a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [15]),
        .Q(\a7/k3a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [16]),
        .Q(\a7/k3a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [17]),
        .Q(\a7/k3a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [18]),
        .Q(\a7/k3a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [19]),
        .Q(\a7/k3a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [1]),
        .Q(\a7/k3a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [20]),
        .Q(\a7/k3a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [21]),
        .Q(\a7/k3a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [22]),
        .Q(\a7/k3a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [23]),
        .Q(\a7/k3a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [24]),
        .Q(\a7/k3a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [25]),
        .Q(\a7/k3a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [26]),
        .Q(\a7/k3a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [27]),
        .Q(\a7/k3a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [28]),
        .Q(\a7/k3a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [29]),
        .Q(\a7/k3a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [2]),
        .Q(\a7/k3a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [30]),
        .Q(\a7/k3a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [31]),
        .Q(\a7/k3a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [3]),
        .Q(\a7/k3a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [4]),
        .Q(\a7/k3a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [5]),
        .Q(\a7/k3a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [6]),
        .Q(\a7/k3a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [7]),
        .Q(\a7/k3a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [8]),
        .Q(\a7/k3a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/k3a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a7/v3 [9]),
        .Q(\a7/k3a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[0]),
        .Q(k7[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[100] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[100]),
        .Q(k7[100]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[101] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[101]),
        .Q(k7[101]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[102] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[102]),
        .Q(k7[102]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[103] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[103]),
        .Q(k7[103]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[104] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[104]),
        .Q(k7[104]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[105] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[105]),
        .Q(k7[105]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[106] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[106]),
        .Q(k7[106]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[107] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[107]),
        .Q(k7[107]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[108] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[108]),
        .Q(k7[108]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[109] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[109]),
        .Q(k7[109]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[10]),
        .Q(k7[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[110] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[110]),
        .Q(k7[110]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[111] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[111]),
        .Q(k7[111]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[112] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[112]),
        .Q(k7[112]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[113] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[113]),
        .Q(k7[113]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[114] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[114]),
        .Q(k7[114]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[115] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[115]),
        .Q(k7[115]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[116] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[116]),
        .Q(k7[116]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[117] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[117]),
        .Q(k7[117]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[118] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[118]),
        .Q(k7[118]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[119] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[119]),
        .Q(k7[119]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[11]),
        .Q(k7[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[120] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[120]),
        .Q(k7[120]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[121] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[121]),
        .Q(k7[121]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[122] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[122]),
        .Q(k7[122]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[123] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[123]),
        .Q(k7[123]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[124] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[124]),
        .Q(k7[124]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[125] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[125]),
        .Q(k7[125]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[126] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[126]),
        .Q(k7[126]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[127] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[127]),
        .Q(k7[127]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[12]),
        .Q(k7[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[13]),
        .Q(k7[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[14]),
        .Q(k7[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[15]),
        .Q(k7[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[16]),
        .Q(k7[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[17]),
        .Q(k7[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[18]),
        .Q(k7[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[19]),
        .Q(k7[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[1]),
        .Q(k7[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[20]),
        .Q(k7[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[21]),
        .Q(k7[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[22]),
        .Q(k7[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[23]),
        .Q(k7[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[24]),
        .Q(k7[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[25]),
        .Q(k7[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[26]),
        .Q(k7[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[27]),
        .Q(k7[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[28]),
        .Q(k7[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[29]),
        .Q(k7[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[2]),
        .Q(k7[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[30]),
        .Q(k7[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[31]),
        .Q(k7[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[32]),
        .Q(k7[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[33]),
        .Q(k7[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[34]),
        .Q(k7[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[35]),
        .Q(k7[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[36]),
        .Q(k7[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[37]),
        .Q(k7[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[38]),
        .Q(k7[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[39]),
        .Q(k7[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[3]),
        .Q(k7[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[40]),
        .Q(k7[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[41]),
        .Q(k7[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[42]),
        .Q(k7[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[43]),
        .Q(k7[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[44]),
        .Q(k7[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[45]),
        .Q(k7[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[46]),
        .Q(k7[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[47]),
        .Q(k7[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[48]),
        .Q(k7[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[49]),
        .Q(k7[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[4]),
        .Q(k7[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[50]),
        .Q(k7[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[51]),
        .Q(k7[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[52]),
        .Q(k7[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[53]),
        .Q(k7[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[54]),
        .Q(k7[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[55]),
        .Q(k7[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[56]),
        .Q(k7[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[57]),
        .Q(k7[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[58]),
        .Q(k7[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[59]),
        .Q(k7[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[5]),
        .Q(k7[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[60]),
        .Q(k7[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[61]),
        .Q(k7[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[62]),
        .Q(k7[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[63]),
        .Q(k7[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[64] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[64]),
        .Q(k7[64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[65] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[65]),
        .Q(k7[65]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[66] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[66]),
        .Q(k7[66]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[67] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[67]),
        .Q(k7[67]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[68] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[68]),
        .Q(k7[68]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[69] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[69]),
        .Q(k7[69]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[6]),
        .Q(k7[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[70] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[70]),
        .Q(k7[70]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[71] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[71]),
        .Q(k7[71]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[72] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[72]),
        .Q(k7[72]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[73] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[73]),
        .Q(k7[73]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[74] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[74]),
        .Q(k7[74]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[75] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[75]),
        .Q(k7[75]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[76] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[76]),
        .Q(k7[76]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[77] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[77]),
        .Q(k7[77]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[78] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[78]),
        .Q(k7[78]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[79] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[79]),
        .Q(k7[79]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[7]),
        .Q(k7[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[80] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[80]),
        .Q(k7[80]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[81] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[81]),
        .Q(k7[81]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[82] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[82]),
        .Q(k7[82]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[83] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[83]),
        .Q(k7[83]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[84] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[84]),
        .Q(k7[84]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[85] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[85]),
        .Q(k7[85]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[86] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[86]),
        .Q(k7[86]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[87] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[87]),
        .Q(k7[87]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[88] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[88]),
        .Q(k7[88]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[89] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[89]),
        .Q(k7[89]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[8]),
        .Q(k7[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[90] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[90]),
        .Q(k7[90]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[91] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[91]),
        .Q(k7[91]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[92] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[92]),
        .Q(k7[92]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[93] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[93]),
        .Q(k7[93]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[94] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[94]),
        .Q(k7[94]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[95] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[95]),
        .Q(k7[95]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[96] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[96]),
        .Q(k7[96]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[97] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[97]),
        .Q(k7[97]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[98] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[98]),
        .Q(k7[98]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[99] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[99]),
        .Q(k7[99]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a7/out_1_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k6b[9]),
        .Q(k7[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_0/S_1/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \a8/S4_0/S_1/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,k7[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,k7[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\a8/S4_0/S_1/out_reg_n_0 ,\a8/S4_0/S_1/out_reg_n_1 ,\a8/S4_0/S_1/out_reg_n_2 ,\a8/S4_0/S_1/out_reg_n_3 ,\a8/S4_0/S_1/out_reg_n_4 ,\a8/S4_0/S_1/out_reg_n_5 ,\a8/S4_0/S_1/out_reg_n_6 ,\a8/S4_0/S_1/out_reg_n_7 ,\a8/k4a [23:16]}),
        .DOBDO({\a8/S4_0/S_1/out_reg_n_16 ,\a8/S4_0/S_1/out_reg_n_17 ,\a8/S4_0/S_1/out_reg_n_18 ,\a8/S4_0/S_1/out_reg_n_19 ,\a8/S4_0/S_1/out_reg_n_20 ,\a8/S4_0/S_1/out_reg_n_21 ,\a8/S4_0/S_1/out_reg_n_22 ,\a8/S4_0/S_1/out_reg_n_23 ,\a8/k4a [31:24]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_0/S_3/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \a8/S4_0/S_3/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,k7[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,k7[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\a8/S4_0/S_3/out_reg_n_0 ,\a8/S4_0/S_3/out_reg_n_1 ,\a8/S4_0/S_3/out_reg_n_2 ,\a8/S4_0/S_3/out_reg_n_3 ,\a8/S4_0/S_3/out_reg_n_4 ,\a8/S4_0/S_3/out_reg_n_5 ,\a8/S4_0/S_3/out_reg_n_6 ,\a8/S4_0/S_3/out_reg_n_7 ,\a8/k4a [7:0]}),
        .DOBDO({\a8/S4_0/S_3/out_reg_n_16 ,\a8/S4_0/S_3/out_reg_n_17 ,\a8/S4_0/S_3/out_reg_n_18 ,\a8/S4_0/S_3/out_reg_n_19 ,\a8/S4_0/S_3/out_reg_n_20 ,\a8/S4_0/S_3/out_reg_n_21 ,\a8/S4_0/S_3/out_reg_n_22 ,\a8/S4_0/S_3/out_reg_n_23 ,\a8/k4a [15:8]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[96]),
        .Q(\a8/k0a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[106]),
        .Q(\a8/k0a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[107]),
        .Q(\a8/k0a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[108]),
        .Q(\a8/k0a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[109]),
        .Q(\a8/k0a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[110]),
        .Q(\a8/k0a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[111]),
        .Q(\a8/k0a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[112]),
        .Q(\a8/k0a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[113]),
        .Q(\a8/k0a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[114]),
        .Q(\a8/k0a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[115]),
        .Q(\a8/k0a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[97]),
        .Q(\a8/k0a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[116]),
        .Q(\a8/k0a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[117]),
        .Q(\a8/k0a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[118]),
        .Q(\a8/k0a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[119]),
        .Q(\a8/k0a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[120]),
        .Q(\a8/k0a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[121]),
        .Q(\a8/k0a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[122]),
        .Q(\a8/k0a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[123]),
        .Q(\a8/k0a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[124]),
        .Q(\a8/k0a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[125]),
        .Q(\a8/k0a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[98]),
        .Q(\a8/k0a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[126]),
        .Q(\a8/k0a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v0 ),
        .Q(\a8/k0a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[99]),
        .Q(\a8/k0a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[100]),
        .Q(\a8/k0a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[101]),
        .Q(\a8/k0a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[102]),
        .Q(\a8/k0a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[103]),
        .Q(\a8/k0a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[104]),
        .Q(\a8/k0a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k0a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7[105]),
        .Q(\a8/k0a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [0]),
        .Q(\a8/k1a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [10]),
        .Q(\a8/k1a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [11]),
        .Q(\a8/k1a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [12]),
        .Q(\a8/k1a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [13]),
        .Q(\a8/k1a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [14]),
        .Q(\a8/k1a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [15]),
        .Q(\a8/k1a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [16]),
        .Q(\a8/k1a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [17]),
        .Q(\a8/k1a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [18]),
        .Q(\a8/k1a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [19]),
        .Q(\a8/k1a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [1]),
        .Q(\a8/k1a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [20]),
        .Q(\a8/k1a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [21]),
        .Q(\a8/k1a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [22]),
        .Q(\a8/k1a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [23]),
        .Q(\a8/k1a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [24]),
        .Q(\a8/k1a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [25]),
        .Q(\a8/k1a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [26]),
        .Q(\a8/k1a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [27]),
        .Q(\a8/k1a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [28]),
        .Q(\a8/k1a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [29]),
        .Q(\a8/k1a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [2]),
        .Q(\a8/k1a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [30]),
        .Q(\a8/k1a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\k1a[31]_i_1__6_n_0 ),
        .Q(\a8/k1a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [3]),
        .Q(\a8/k1a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [4]),
        .Q(\a8/k1a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [5]),
        .Q(\a8/k1a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [6]),
        .Q(\a8/k1a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [7]),
        .Q(\a8/k1a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [8]),
        .Q(\a8/k1a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k1a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v1 [9]),
        .Q(\a8/k1a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [0]),
        .Q(\a8/k2a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [10]),
        .Q(\a8/k2a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [11]),
        .Q(\a8/k2a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [12]),
        .Q(\a8/k2a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [13]),
        .Q(\a8/k2a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [14]),
        .Q(\a8/k2a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [15]),
        .Q(\a8/k2a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [16]),
        .Q(\a8/k2a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [17]),
        .Q(\a8/k2a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [18]),
        .Q(\a8/k2a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [19]),
        .Q(\a8/k2a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [1]),
        .Q(\a8/k2a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [20]),
        .Q(\a8/k2a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [21]),
        .Q(\a8/k2a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [22]),
        .Q(\a8/k2a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [23]),
        .Q(\a8/k2a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [24]),
        .Q(\a8/k2a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [25]),
        .Q(\a8/k2a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [26]),
        .Q(\a8/k2a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [27]),
        .Q(\a8/k2a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [28]),
        .Q(\a8/k2a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [29]),
        .Q(\a8/k2a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [2]),
        .Q(\a8/k2a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [30]),
        .Q(\a8/k2a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [31]),
        .Q(\a8/k2a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [3]),
        .Q(\a8/k2a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [4]),
        .Q(\a8/k2a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [5]),
        .Q(\a8/k2a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [6]),
        .Q(\a8/k2a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [7]),
        .Q(\a8/k2a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [8]),
        .Q(\a8/k2a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k2a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v2 [9]),
        .Q(\a8/k2a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [0]),
        .Q(\a8/k3a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [10]),
        .Q(\a8/k3a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [11]),
        .Q(\a8/k3a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [12]),
        .Q(\a8/k3a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [13]),
        .Q(\a8/k3a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [14]),
        .Q(\a8/k3a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [15]),
        .Q(\a8/k3a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [16]),
        .Q(\a8/k3a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [17]),
        .Q(\a8/k3a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [18]),
        .Q(\a8/k3a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [19]),
        .Q(\a8/k3a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [1]),
        .Q(\a8/k3a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [20]),
        .Q(\a8/k3a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [21]),
        .Q(\a8/k3a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [22]),
        .Q(\a8/k3a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [23]),
        .Q(\a8/k3a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [24]),
        .Q(\a8/k3a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [25]),
        .Q(\a8/k3a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [26]),
        .Q(\a8/k3a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [27]),
        .Q(\a8/k3a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [28]),
        .Q(\a8/k3a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [29]),
        .Q(\a8/k3a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [2]),
        .Q(\a8/k3a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [30]),
        .Q(\a8/k3a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [31]),
        .Q(\a8/k3a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [3]),
        .Q(\a8/k3a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [4]),
        .Q(\a8/k3a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [5]),
        .Q(\a8/k3a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [6]),
        .Q(\a8/k3a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [7]),
        .Q(\a8/k3a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [8]),
        .Q(\a8/k3a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/k3a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a8/v3 [9]),
        .Q(\a8/k3a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[0]),
        .Q(k8[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[100] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[100]),
        .Q(k8[100]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[101] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[101]),
        .Q(k8[101]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[102] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[102]),
        .Q(k8[102]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[103] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[103]),
        .Q(k8[103]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[104] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[104]),
        .Q(k8[104]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[105] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[105]),
        .Q(k8[105]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[106] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[106]),
        .Q(k8[106]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[107] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[107]),
        .Q(k8[107]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[108] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[108]),
        .Q(k8[108]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[109] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[109]),
        .Q(k8[109]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[10]),
        .Q(k8[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[110] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[110]),
        .Q(k8[110]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[111] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[111]),
        .Q(k8[111]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[112] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[112]),
        .Q(k8[112]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[113] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[113]),
        .Q(k8[113]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[114] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[114]),
        .Q(k8[114]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[115] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[115]),
        .Q(k8[115]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[116] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[116]),
        .Q(k8[116]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[117] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[117]),
        .Q(k8[117]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[118] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[118]),
        .Q(k8[118]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[119] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[119]),
        .Q(k8[119]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[11]),
        .Q(k8[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[120] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[120]),
        .Q(k8[120]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[121] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[121]),
        .Q(k8[121]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[122] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[122]),
        .Q(k8[122]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[123] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[123]),
        .Q(k8[123]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[124] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[124]),
        .Q(k8[124]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[125] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[125]),
        .Q(k8[125]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[126] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[126]),
        .Q(k8[126]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[127] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[127]),
        .Q(k8[127]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[12]),
        .Q(k8[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[13]),
        .Q(k8[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[14]),
        .Q(k8[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[15]),
        .Q(k8[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[16]),
        .Q(k8[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[17]),
        .Q(k8[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[18]),
        .Q(k8[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[19]),
        .Q(k8[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[1]),
        .Q(k8[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[20]),
        .Q(k8[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[21]),
        .Q(k8[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[22]),
        .Q(k8[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[23]),
        .Q(k8[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[24]),
        .Q(k8[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[25]),
        .Q(k8[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[26]),
        .Q(k8[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[27]),
        .Q(k8[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[28]),
        .Q(k8[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[29]),
        .Q(k8[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[2]),
        .Q(k8[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[30]),
        .Q(k8[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[31]),
        .Q(k8[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[32]),
        .Q(k8[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[33]),
        .Q(k8[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[34]),
        .Q(k8[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[35]),
        .Q(k8[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[36]),
        .Q(k8[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[37]),
        .Q(k8[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[38]),
        .Q(k8[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[39]),
        .Q(k8[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[3]),
        .Q(k8[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[40]),
        .Q(k8[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[41]),
        .Q(k8[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[42]),
        .Q(k8[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[43]),
        .Q(k8[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[44]),
        .Q(k8[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[45]),
        .Q(k8[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[46]),
        .Q(k8[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[47]),
        .Q(k8[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[48]),
        .Q(k8[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[49]),
        .Q(k8[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[4]),
        .Q(k8[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[50]),
        .Q(k8[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[51]),
        .Q(k8[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[52]),
        .Q(k8[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[53]),
        .Q(k8[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[54]),
        .Q(k8[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[55]),
        .Q(k8[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[56]),
        .Q(k8[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[57]),
        .Q(k8[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[58]),
        .Q(k8[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[59]),
        .Q(k8[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[5]),
        .Q(k8[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[60]),
        .Q(k8[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[61]),
        .Q(k8[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[62]),
        .Q(k8[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[63]),
        .Q(k8[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[64] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[64]),
        .Q(k8[64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[65] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[65]),
        .Q(k8[65]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[66] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[66]),
        .Q(k8[66]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[67] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[67]),
        .Q(k8[67]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[68] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[68]),
        .Q(k8[68]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[69] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[69]),
        .Q(k8[69]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[6]),
        .Q(k8[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[70] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[70]),
        .Q(k8[70]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[71] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[71]),
        .Q(k8[71]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[72] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[72]),
        .Q(k8[72]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[73] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[73]),
        .Q(k8[73]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[74] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[74]),
        .Q(k8[74]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[75] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[75]),
        .Q(k8[75]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[76] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[76]),
        .Q(k8[76]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[77] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[77]),
        .Q(k8[77]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[78] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[78]),
        .Q(k8[78]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[79] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[79]),
        .Q(k8[79]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[7]),
        .Q(k8[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[80] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[80]),
        .Q(k8[80]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[81] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[81]),
        .Q(k8[81]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[82] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[82]),
        .Q(k8[82]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[83] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[83]),
        .Q(k8[83]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[84] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[84]),
        .Q(k8[84]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[85] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[85]),
        .Q(k8[85]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[86] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[86]),
        .Q(k8[86]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[87] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[87]),
        .Q(k8[87]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[88] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[88]),
        .Q(k8[88]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[89] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[89]),
        .Q(k8[89]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[8]),
        .Q(k8[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[90] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[90]),
        .Q(k8[90]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[91] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[91]),
        .Q(k8[91]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[92] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[92]),
        .Q(k8[92]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[93] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[93]),
        .Q(k8[93]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[94] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[94]),
        .Q(k8[94]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[95] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[95]),
        .Q(k8[95]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[96] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[96]),
        .Q(k8[96]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[97] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[97]),
        .Q(k8[97]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[98] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[98]),
        .Q(k8[98]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[99] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[99]),
        .Q(k8[99]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a8/out_1_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k7b[9]),
        .Q(k8[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_0/S_1/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \a9/S4_0/S_1/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,k8[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,k8[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\a9/S4_0/S_1/out_reg_n_0 ,\a9/S4_0/S_1/out_reg_n_1 ,\a9/S4_0/S_1/out_reg_n_2 ,\a9/S4_0/S_1/out_reg_n_3 ,\a9/S4_0/S_1/out_reg_n_4 ,\a9/S4_0/S_1/out_reg_n_5 ,\a9/S4_0/S_1/out_reg_n_6 ,\a9/S4_0/S_1/out_reg_n_7 ,\a9/k4a [23:16]}),
        .DOBDO({\a9/S4_0/S_1/out_reg_n_16 ,\a9/S4_0/S_1/out_reg_n_17 ,\a9/S4_0/S_1/out_reg_n_18 ,\a9/S4_0/S_1/out_reg_n_19 ,\a9/S4_0/S_1/out_reg_n_20 ,\a9/S4_0/S_1/out_reg_n_21 ,\a9/S4_0/S_1/out_reg_n_22 ,\a9/S4_0/S_1/out_reg_n_23 ,\a9/k4a [31:24]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_0/S_3/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \a9/S4_0/S_3/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,k8[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,k8[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\a9/S4_0/S_3/out_reg_n_0 ,\a9/S4_0/S_3/out_reg_n_1 ,\a9/S4_0/S_3/out_reg_n_2 ,\a9/S4_0/S_3/out_reg_n_3 ,\a9/S4_0/S_3/out_reg_n_4 ,\a9/S4_0/S_3/out_reg_n_5 ,\a9/S4_0/S_3/out_reg_n_6 ,\a9/S4_0/S_3/out_reg_n_7 ,\a9/k4a [7:0]}),
        .DOBDO({\a9/S4_0/S_3/out_reg_n_16 ,\a9/S4_0/S_3/out_reg_n_17 ,\a9/S4_0/S_3/out_reg_n_18 ,\a9/S4_0/S_3/out_reg_n_19 ,\a9/S4_0/S_3/out_reg_n_20 ,\a9/S4_0/S_3/out_reg_n_21 ,\a9/S4_0/S_3/out_reg_n_22 ,\a9/S4_0/S_3/out_reg_n_23 ,\a9/k4a [15:8]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[96]),
        .Q(\a9/k0a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[106]),
        .Q(\a9/k0a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[107]),
        .Q(\a9/k0a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[108]),
        .Q(\a9/k0a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[109]),
        .Q(\a9/k0a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[110]),
        .Q(\a9/k0a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[111]),
        .Q(\a9/k0a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[112]),
        .Q(\a9/k0a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[113]),
        .Q(\a9/k0a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[114]),
        .Q(\a9/k0a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[115]),
        .Q(\a9/k0a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[97]),
        .Q(\a9/k0a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[116]),
        .Q(\a9/k0a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[117]),
        .Q(\a9/k0a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[118]),
        .Q(\a9/k0a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[119]),
        .Q(\a9/k0a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v0 [24]),
        .Q(\a9/k0a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v0 [25]),
        .Q(\a9/k0a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[122]),
        .Q(\a9/k0a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v0 [27]),
        .Q(\a9/k0a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v0 [28]),
        .Q(\a9/k0a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[125]),
        .Q(\a9/k0a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[98]),
        .Q(\a9/k0a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[126]),
        .Q(\a9/k0a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[127]),
        .Q(\a9/k0a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[99]),
        .Q(\a9/k0a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[100]),
        .Q(\a9/k0a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[101]),
        .Q(\a9/k0a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[102]),
        .Q(\a9/k0a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[103]),
        .Q(\a9/k0a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[104]),
        .Q(\a9/k0a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k0a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8[105]),
        .Q(\a9/k0a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [0]),
        .Q(\a9/k1a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [10]),
        .Q(\a9/k1a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [11]),
        .Q(\a9/k1a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [12]),
        .Q(\a9/k1a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [13]),
        .Q(\a9/k1a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [14]),
        .Q(\a9/k1a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [15]),
        .Q(\a9/k1a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [16]),
        .Q(\a9/k1a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [17]),
        .Q(\a9/k1a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [18]),
        .Q(\a9/k1a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [19]),
        .Q(\a9/k1a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [1]),
        .Q(\a9/k1a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [20]),
        .Q(\a9/k1a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [21]),
        .Q(\a9/k1a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [22]),
        .Q(\a9/k1a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [23]),
        .Q(\a9/k1a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k1a),
        .Q(\a9/k1a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\k1a[25]_i_1__7_n_0 ),
        .Q(\a9/k1a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [26]),
        .Q(\a9/k1a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\k1a[27]_i_1__7_n_0 ),
        .Q(\a9/k1a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\k1a[28]_i_1__7_n_0 ),
        .Q(\a9/k1a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [29]),
        .Q(\a9/k1a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [2]),
        .Q(\a9/k1a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [30]),
        .Q(\a9/k1a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [31]),
        .Q(\a9/k1a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [3]),
        .Q(\a9/k1a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [4]),
        .Q(\a9/k1a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [5]),
        .Q(\a9/k1a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [6]),
        .Q(\a9/k1a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [7]),
        .Q(\a9/k1a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [8]),
        .Q(\a9/k1a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k1a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v1 [9]),
        .Q(\a9/k1a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [0]),
        .Q(\a9/k2a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [10]),
        .Q(\a9/k2a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [11]),
        .Q(\a9/k2a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [12]),
        .Q(\a9/k2a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [13]),
        .Q(\a9/k2a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [14]),
        .Q(\a9/k2a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [15]),
        .Q(\a9/k2a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [16]),
        .Q(\a9/k2a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [17]),
        .Q(\a9/k2a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [18]),
        .Q(\a9/k2a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [19]),
        .Q(\a9/k2a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [1]),
        .Q(\a9/k2a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [20]),
        .Q(\a9/k2a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [21]),
        .Q(\a9/k2a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [22]),
        .Q(\a9/k2a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [23]),
        .Q(\a9/k2a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [24]),
        .Q(\a9/k2a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [25]),
        .Q(\a9/k2a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [26]),
        .Q(\a9/k2a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [27]),
        .Q(\a9/k2a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [28]),
        .Q(\a9/k2a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [29]),
        .Q(\a9/k2a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [2]),
        .Q(\a9/k2a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [30]),
        .Q(\a9/k2a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [31]),
        .Q(\a9/k2a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [3]),
        .Q(\a9/k2a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [4]),
        .Q(\a9/k2a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [5]),
        .Q(\a9/k2a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [6]),
        .Q(\a9/k2a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [7]),
        .Q(\a9/k2a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [8]),
        .Q(\a9/k2a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k2a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v2 [9]),
        .Q(\a9/k2a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [0]),
        .Q(\a9/k3a [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [10]),
        .Q(\a9/k3a [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [11]),
        .Q(\a9/k3a [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [12]),
        .Q(\a9/k3a [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [13]),
        .Q(\a9/k3a [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [14]),
        .Q(\a9/k3a [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [15]),
        .Q(\a9/k3a [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [16]),
        .Q(\a9/k3a [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [17]),
        .Q(\a9/k3a [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [18]),
        .Q(\a9/k3a [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [19]),
        .Q(\a9/k3a [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [1]),
        .Q(\a9/k3a [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [20]),
        .Q(\a9/k3a [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [21]),
        .Q(\a9/k3a [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [22]),
        .Q(\a9/k3a [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [23]),
        .Q(\a9/k3a [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [24]),
        .Q(\a9/k3a [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [25]),
        .Q(\a9/k3a [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [26]),
        .Q(\a9/k3a [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [27]),
        .Q(\a9/k3a [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [28]),
        .Q(\a9/k3a [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [29]),
        .Q(\a9/k3a [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [2]),
        .Q(\a9/k3a [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [30]),
        .Q(\a9/k3a [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [31]),
        .Q(\a9/k3a [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [3]),
        .Q(\a9/k3a [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [4]),
        .Q(\a9/k3a [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [5]),
        .Q(\a9/k3a [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [6]),
        .Q(\a9/k3a [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [7]),
        .Q(\a9/k3a [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [8]),
        .Q(\a9/k3a [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/k3a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\a9/v3 [9]),
        .Q(\a9/k3a [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[0]),
        .Q(k9[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[100] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[100]),
        .Q(k9[100]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[101] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[101]),
        .Q(k9[101]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[102] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[102]),
        .Q(k9[102]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[103] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[103]),
        .Q(k9[103]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[104] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[104]),
        .Q(k9[104]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[105] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[105]),
        .Q(k9[105]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[106] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[106]),
        .Q(k9[106]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[107] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[107]),
        .Q(k9[107]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[108] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[108]),
        .Q(k9[108]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[109] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[109]),
        .Q(k9[109]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[10]),
        .Q(k9[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[110] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[110]),
        .Q(k9[110]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[111] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[111]),
        .Q(k9[111]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[112] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[112]),
        .Q(k9[112]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[113] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[113]),
        .Q(k9[113]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[114] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[114]),
        .Q(k9[114]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[115] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[115]),
        .Q(k9[115]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[116] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[116]),
        .Q(k9[116]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[117] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[117]),
        .Q(k9[117]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[118] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[118]),
        .Q(k9[118]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[119] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[119]),
        .Q(k9[119]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[11]),
        .Q(k9[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[120] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[120]),
        .Q(k9[120]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[121] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[121]),
        .Q(k9[121]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[122] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[122]),
        .Q(k9[122]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[123] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[123]),
        .Q(k9[123]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[124] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[124]),
        .Q(k9[124]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[125] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[125]),
        .Q(k9[125]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[126] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[126]),
        .Q(k9[126]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[127] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[127]),
        .Q(k9[127]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[12]),
        .Q(k9[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[13]),
        .Q(k9[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[14]),
        .Q(k9[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[15]),
        .Q(k9[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[16]),
        .Q(k9[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[17]),
        .Q(k9[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[18]),
        .Q(k9[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[19]),
        .Q(k9[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[1]),
        .Q(k9[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[20]),
        .Q(k9[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[21]),
        .Q(k9[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[22]),
        .Q(k9[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[23]),
        .Q(k9[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[24]),
        .Q(k9[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[25]),
        .Q(k9[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[26]),
        .Q(k9[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[27]),
        .Q(k9[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[28]),
        .Q(k9[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[29]),
        .Q(k9[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[2]),
        .Q(k9[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[30]),
        .Q(k9[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[31]),
        .Q(k9[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[32]),
        .Q(k9[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[33]),
        .Q(k9[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[34]),
        .Q(k9[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[35]),
        .Q(k9[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[36]),
        .Q(k9[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[37]),
        .Q(k9[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[38]),
        .Q(k9[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[39]),
        .Q(k9[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[3]),
        .Q(k9[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[40]),
        .Q(k9[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[41]),
        .Q(k9[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[42]),
        .Q(k9[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[43]),
        .Q(k9[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[44]),
        .Q(k9[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[45]),
        .Q(k9[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[46]),
        .Q(k9[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[47]),
        .Q(k9[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[48]),
        .Q(k9[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[49]),
        .Q(k9[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[4]),
        .Q(k9[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[50]),
        .Q(k9[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[51]),
        .Q(k9[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[52]),
        .Q(k9[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[53]),
        .Q(k9[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[54]),
        .Q(k9[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[55]),
        .Q(k9[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[56]),
        .Q(k9[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[57]),
        .Q(k9[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[58]),
        .Q(k9[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[59]),
        .Q(k9[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[5]),
        .Q(k9[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[60]),
        .Q(k9[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[61]),
        .Q(k9[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[62]),
        .Q(k9[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[63]),
        .Q(k9[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[64] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[64]),
        .Q(k9[64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[65] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[65]),
        .Q(k9[65]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[66] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[66]),
        .Q(k9[66]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[67] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[67]),
        .Q(k9[67]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[68] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[68]),
        .Q(k9[68]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[69] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[69]),
        .Q(k9[69]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[6]),
        .Q(k9[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[70] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[70]),
        .Q(k9[70]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[71] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[71]),
        .Q(k9[71]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[72] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[72]),
        .Q(k9[72]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[73] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[73]),
        .Q(k9[73]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[74] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[74]),
        .Q(k9[74]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[75] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[75]),
        .Q(k9[75]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[76] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[76]),
        .Q(k9[76]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[77] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[77]),
        .Q(k9[77]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[78] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[78]),
        .Q(k9[78]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[79] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[79]),
        .Q(k9[79]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[7]),
        .Q(k9[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[80] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[80]),
        .Q(k9[80]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[81] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[81]),
        .Q(k9[81]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[82] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[82]),
        .Q(k9[82]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[83] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[83]),
        .Q(k9[83]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[84] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[84]),
        .Q(k9[84]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[85] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[85]),
        .Q(k9[85]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[86] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[86]),
        .Q(k9[86]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[87] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[87]),
        .Q(k9[87]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[88] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[88]),
        .Q(k9[88]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[89] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[89]),
        .Q(k9[89]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[8]),
        .Q(k9[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[90] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[90]),
        .Q(k9[90]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[91] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[91]),
        .Q(k9[91]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[92] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[92]),
        .Q(k9[92]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[93] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[93]),
        .Q(k9[93]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[94] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[94]),
        .Q(k9[94]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[95] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[95]),
        .Q(k9[95]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[96] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[96]),
        .Q(k9[96]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[97] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[97]),
        .Q(k9[97]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[98] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[98]),
        .Q(k9[98]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[99] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[99]),
        .Q(k9[99]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \a9/out_1_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(k8b[9]),
        .Q(k9[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[0]),
        .Q(k0[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[100] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[100]),
        .Q(k0[100]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[101] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[101]),
        .Q(k0[101]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[102] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[102]),
        .Q(k0[102]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[103] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[103]),
        .Q(k0[103]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[104] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[104]),
        .Q(k0[104]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[105] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[105]),
        .Q(k0[105]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[106] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[106]),
        .Q(k0[106]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[107] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[107]),
        .Q(k0[107]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[108] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[108]),
        .Q(k0[108]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[109] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[109]),
        .Q(k0[109]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[10]),
        .Q(k0[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[110] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[110]),
        .Q(k0[110]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[111] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[111]),
        .Q(k0[111]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[112] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[112]),
        .Q(k0[112]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[113] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[113]),
        .Q(k0[113]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[114] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[114]),
        .Q(k0[114]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[115] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[115]),
        .Q(k0[115]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[116] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[116]),
        .Q(k0[116]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[117] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[117]),
        .Q(k0[117]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[118] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[118]),
        .Q(k0[118]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[119] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[119]),
        .Q(k0[119]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[11]),
        .Q(k0[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[120] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[120]),
        .Q(k0[120]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[121] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[121]),
        .Q(k0[121]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[122] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[122]),
        .Q(k0[122]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[123] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[123]),
        .Q(k0[123]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[124] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[124]),
        .Q(k0[124]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[125] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[125]),
        .Q(k0[125]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[126] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[126]),
        .Q(k0[126]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[127] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[127]),
        .Q(k0[127]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[12]),
        .Q(k0[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[13]),
        .Q(k0[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[14]),
        .Q(k0[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[15]),
        .Q(k0[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[16]),
        .Q(k0[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[17]),
        .Q(k0[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[18]),
        .Q(k0[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[19]),
        .Q(k0[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[1]),
        .Q(k0[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[20]),
        .Q(k0[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[21]),
        .Q(k0[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[22]),
        .Q(k0[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[23]),
        .Q(k0[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[24]),
        .Q(k0[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[25]),
        .Q(k0[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[26]),
        .Q(k0[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[27]),
        .Q(k0[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[28]),
        .Q(k0[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[29]),
        .Q(k0[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[2]),
        .Q(k0[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[30]),
        .Q(k0[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[31]),
        .Q(k0[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[32]),
        .Q(k0[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[33]),
        .Q(k0[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[34]),
        .Q(k0[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[35]),
        .Q(k0[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[36]),
        .Q(k0[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[37]),
        .Q(k0[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[38]),
        .Q(k0[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[39]),
        .Q(k0[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[3]),
        .Q(k0[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[40]),
        .Q(k0[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[41]),
        .Q(k0[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[42]),
        .Q(k0[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[43]),
        .Q(k0[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[44]),
        .Q(k0[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[45]),
        .Q(k0[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[46]),
        .Q(k0[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[47]),
        .Q(k0[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[48]),
        .Q(k0[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[49]),
        .Q(k0[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[4]),
        .Q(k0[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[50]),
        .Q(k0[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[51]),
        .Q(k0[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[52]),
        .Q(k0[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[53]),
        .Q(k0[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[54]),
        .Q(k0[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[55]),
        .Q(k0[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[56]),
        .Q(k0[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[57]),
        .Q(k0[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[58]),
        .Q(k0[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[59]),
        .Q(k0[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[5]),
        .Q(k0[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[60]),
        .Q(k0[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[61]),
        .Q(k0[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[62]),
        .Q(k0[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[63]),
        .Q(k0[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[64] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[64]),
        .Q(k0[64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[65] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[65]),
        .Q(k0[65]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[66] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[66]),
        .Q(k0[66]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[67] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[67]),
        .Q(k0[67]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[68] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[68]),
        .Q(k0[68]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[69] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[69]),
        .Q(k0[69]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[6]),
        .Q(k0[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[70] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[70]),
        .Q(k0[70]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[71] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[71]),
        .Q(k0[71]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[72] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[72]),
        .Q(k0[72]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[73] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[73]),
        .Q(k0[73]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[74] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[74]),
        .Q(k0[74]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[75] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[75]),
        .Q(k0[75]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[76] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[76]),
        .Q(k0[76]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[77] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[77]),
        .Q(k0[77]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[78] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[78]),
        .Q(k0[78]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[79] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[79]),
        .Q(k0[79]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[7]),
        .Q(k0[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[80] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[80]),
        .Q(k0[80]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[81] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[81]),
        .Q(k0[81]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[82] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[82]),
        .Q(k0[82]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[83] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[83]),
        .Q(k0[83]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[84] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[84]),
        .Q(k0[84]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[85] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[85]),
        .Q(k0[85]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[86] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[86]),
        .Q(k0[86]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[87] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[87]),
        .Q(k0[87]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[88] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[88]),
        .Q(k0[88]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[89] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[89]),
        .Q(k0[89]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[8]),
        .Q(k0[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[90] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[90]),
        .Q(k0[90]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[91] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[91]),
        .Q(k0[91]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[92] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[92]),
        .Q(k0[92]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[93] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[93]),
        .Q(k0[93]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[94] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[94]),
        .Q(k0[94]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[95] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[95]),
        .Q(k0[95]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[96] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[96]),
        .Q(k0[96]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[97] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[97]),
        .Q(k0[97]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[98] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[98]),
        .Q(k0[98]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[99] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[99]),
        .Q(k0[99]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \k0_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key[9]),
        .Q(k0[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair879" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \k0a[24]_i_1 
       (.I0(k0[120]),
        .O(\a1/v0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair451" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \k0a[24]_i_1__0 
       (.I0(k8[120]),
        .O(\a9/v0 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair814" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \k0a[25]_i_1 
       (.I0(k1[121]),
        .O(\a2/v0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair450" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \k0a[25]_i_1__0 
       (.I0(k8[121]),
        .O(\a9/v0 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair487" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \k0a[25]_i_1__1 
       (.I0(k9[121]),
        .O(\a10/v0 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair749" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \k0a[26]_i_1 
       (.I0(k2[122]),
        .O(\a3/v0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair486" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \k0a[26]_i_1__0 
       (.I0(k9[122]),
        .O(\a10/v0 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair684" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \k0a[27]_i_1 
       (.I0(k3[123]),
        .O(\a4/v0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair449" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \k0a[27]_i_1__0 
       (.I0(k8[123]),
        .O(\a9/v0 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair618" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \k0a[28]_i_1 
       (.I0(k4[124]),
        .O(\a5/v0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair448" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \k0a[28]_i_1__0 
       (.I0(k8[124]),
        .O(\a9/v0 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair485" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \k0a[28]_i_1__1 
       (.I0(k9[124]),
        .O(\a10/v0 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair553" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \k0a[29]_i_1 
       (.I0(k5[125]),
        .O(\a6/v0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair484" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \k0a[29]_i_1__0 
       (.I0(k9[125]),
        .O(\a10/v0 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair488" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \k0a[30]_i_1 
       (.I0(k6[126]),
        .O(\a7/v0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair945" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \k0a[31]_i_1 
       (.I0(k7[127]),
        .O(\a8/v0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[0]_i_1 
       (.I0(k0[96]),
        .I1(k0[64]),
        .O(\a1/v1 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[0]_i_1__0 
       (.I0(k1[96]),
        .I1(k1[64]),
        .O(\a2/v1 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[0]_i_1__1 
       (.I0(k2[96]),
        .I1(k2[64]),
        .O(\a3/v1 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[0]_i_1__2 
       (.I0(k3[96]),
        .I1(k3[64]),
        .O(\a4/v1 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[0]_i_1__3 
       (.I0(k4[96]),
        .I1(k4[64]),
        .O(\a5/v1 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[0]_i_1__4 
       (.I0(k5[96]),
        .I1(k5[64]),
        .O(\a6/v1 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[0]_i_1__5 
       (.I0(k6[96]),
        .I1(k6[64]),
        .O(\a7/v1 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[0]_i_1__6 
       (.I0(k7[96]),
        .I1(k7[64]),
        .O(\a8/v1 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[0]_i_1__7 
       (.I0(k8[96]),
        .I1(k8[64]),
        .O(\a9/v1 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[0]_i_1__8 
       (.I0(k9[96]),
        .I1(k9[64]),
        .O(\a10/v1 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[10]_i_1 
       (.I0(k0[106]),
        .I1(k0[74]),
        .O(\a1/v1 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[10]_i_1__0 
       (.I0(k1[106]),
        .I1(k1[74]),
        .O(\a2/v1 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[10]_i_1__1 
       (.I0(k2[106]),
        .I1(k2[74]),
        .O(\a3/v1 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[10]_i_1__2 
       (.I0(k3[106]),
        .I1(k3[74]),
        .O(\a4/v1 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[10]_i_1__3 
       (.I0(k4[106]),
        .I1(k4[74]),
        .O(\a5/v1 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[10]_i_1__4 
       (.I0(k5[106]),
        .I1(k5[74]),
        .O(\a6/v1 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[10]_i_1__5 
       (.I0(k6[106]),
        .I1(k6[74]),
        .O(\a7/v1 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[10]_i_1__6 
       (.I0(k7[106]),
        .I1(k7[74]),
        .O(\a8/v1 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[10]_i_1__7 
       (.I0(k8[106]),
        .I1(k8[74]),
        .O(\a9/v1 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[10]_i_1__8 
       (.I0(k9[106]),
        .I1(k9[74]),
        .O(\a10/v1 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[11]_i_1 
       (.I0(k0[107]),
        .I1(k0[75]),
        .O(\a1/v1 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[11]_i_1__0 
       (.I0(k1[107]),
        .I1(k1[75]),
        .O(\a2/v1 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[11]_i_1__1 
       (.I0(k2[107]),
        .I1(k2[75]),
        .O(\a3/v1 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[11]_i_1__2 
       (.I0(k3[107]),
        .I1(k3[75]),
        .O(\a4/v1 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[11]_i_1__3 
       (.I0(k4[107]),
        .I1(k4[75]),
        .O(\a5/v1 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[11]_i_1__4 
       (.I0(k5[107]),
        .I1(k5[75]),
        .O(\a6/v1 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[11]_i_1__5 
       (.I0(k6[107]),
        .I1(k6[75]),
        .O(\a7/v1 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[11]_i_1__6 
       (.I0(k7[107]),
        .I1(k7[75]),
        .O(\a8/v1 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[11]_i_1__7 
       (.I0(k8[107]),
        .I1(k8[75]),
        .O(\a9/v1 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[11]_i_1__8 
       (.I0(k9[107]),
        .I1(k9[75]),
        .O(\a10/v1 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[12]_i_1 
       (.I0(k0[108]),
        .I1(k0[76]),
        .O(\a1/v1 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[12]_i_1__0 
       (.I0(k1[108]),
        .I1(k1[76]),
        .O(\a2/v1 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[12]_i_1__1 
       (.I0(k2[108]),
        .I1(k2[76]),
        .O(\a3/v1 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[12]_i_1__2 
       (.I0(k3[108]),
        .I1(k3[76]),
        .O(\a4/v1 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[12]_i_1__3 
       (.I0(k4[108]),
        .I1(k4[76]),
        .O(\a5/v1 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[12]_i_1__4 
       (.I0(k5[108]),
        .I1(k5[76]),
        .O(\a6/v1 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[12]_i_1__5 
       (.I0(k6[108]),
        .I1(k6[76]),
        .O(\a7/v1 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[12]_i_1__6 
       (.I0(k7[108]),
        .I1(k7[76]),
        .O(\a8/v1 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[12]_i_1__7 
       (.I0(k8[108]),
        .I1(k8[76]),
        .O(\a9/v1 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[12]_i_1__8 
       (.I0(k9[108]),
        .I1(k9[76]),
        .O(\a10/v1 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[13]_i_1 
       (.I0(k0[109]),
        .I1(k0[77]),
        .O(\a1/v1 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[13]_i_1__0 
       (.I0(k1[109]),
        .I1(k1[77]),
        .O(\a2/v1 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[13]_i_1__1 
       (.I0(k2[109]),
        .I1(k2[77]),
        .O(\a3/v1 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[13]_i_1__2 
       (.I0(k3[109]),
        .I1(k3[77]),
        .O(\a4/v1 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[13]_i_1__3 
       (.I0(k4[109]),
        .I1(k4[77]),
        .O(\a5/v1 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[13]_i_1__4 
       (.I0(k5[109]),
        .I1(k5[77]),
        .O(\a6/v1 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[13]_i_1__5 
       (.I0(k6[109]),
        .I1(k6[77]),
        .O(\a7/v1 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[13]_i_1__6 
       (.I0(k7[109]),
        .I1(k7[77]),
        .O(\a8/v1 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[13]_i_1__7 
       (.I0(k8[109]),
        .I1(k8[77]),
        .O(\a9/v1 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[13]_i_1__8 
       (.I0(k9[109]),
        .I1(k9[77]),
        .O(\a10/v1 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[14]_i_1 
       (.I0(k0[110]),
        .I1(k0[78]),
        .O(\a1/v1 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[14]_i_1__0 
       (.I0(k1[110]),
        .I1(k1[78]),
        .O(\a2/v1 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[14]_i_1__1 
       (.I0(k2[110]),
        .I1(k2[78]),
        .O(\a3/v1 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[14]_i_1__2 
       (.I0(k3[110]),
        .I1(k3[78]),
        .O(\a4/v1 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[14]_i_1__3 
       (.I0(k4[110]),
        .I1(k4[78]),
        .O(\a5/v1 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[14]_i_1__4 
       (.I0(k5[110]),
        .I1(k5[78]),
        .O(\a6/v1 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[14]_i_1__5 
       (.I0(k6[110]),
        .I1(k6[78]),
        .O(\a7/v1 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[14]_i_1__6 
       (.I0(k7[110]),
        .I1(k7[78]),
        .O(\a8/v1 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[14]_i_1__7 
       (.I0(k8[110]),
        .I1(k8[78]),
        .O(\a9/v1 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[14]_i_1__8 
       (.I0(k9[110]),
        .I1(k9[78]),
        .O(\a10/v1 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[15]_i_1 
       (.I0(k0[111]),
        .I1(k0[79]),
        .O(\a1/v1 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[15]_i_1__0 
       (.I0(k1[111]),
        .I1(k1[79]),
        .O(\a2/v1 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[15]_i_1__1 
       (.I0(k2[111]),
        .I1(k2[79]),
        .O(\a3/v1 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[15]_i_1__2 
       (.I0(k3[111]),
        .I1(k3[79]),
        .O(\a4/v1 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[15]_i_1__3 
       (.I0(k4[111]),
        .I1(k4[79]),
        .O(\a5/v1 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[15]_i_1__4 
       (.I0(k5[111]),
        .I1(k5[79]),
        .O(\a6/v1 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[15]_i_1__5 
       (.I0(k6[111]),
        .I1(k6[79]),
        .O(\a7/v1 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[15]_i_1__6 
       (.I0(k7[111]),
        .I1(k7[79]),
        .O(\a8/v1 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[15]_i_1__7 
       (.I0(k8[111]),
        .I1(k8[79]),
        .O(\a9/v1 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[15]_i_1__8 
       (.I0(k9[111]),
        .I1(k9[79]),
        .O(\a10/v1 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[16]_i_1 
       (.I0(k0[112]),
        .I1(k0[80]),
        .O(\a1/v1 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[16]_i_1__0 
       (.I0(k1[112]),
        .I1(k1[80]),
        .O(\a2/v1 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[16]_i_1__1 
       (.I0(k2[112]),
        .I1(k2[80]),
        .O(\a3/v1 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[16]_i_1__2 
       (.I0(k3[112]),
        .I1(k3[80]),
        .O(\a4/v1 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[16]_i_1__3 
       (.I0(k4[112]),
        .I1(k4[80]),
        .O(\a5/v1 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[16]_i_1__4 
       (.I0(k5[112]),
        .I1(k5[80]),
        .O(\a6/v1 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[16]_i_1__5 
       (.I0(k6[112]),
        .I1(k6[80]),
        .O(\a7/v1 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[16]_i_1__6 
       (.I0(k7[112]),
        .I1(k7[80]),
        .O(\a8/v1 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[16]_i_1__7 
       (.I0(k8[112]),
        .I1(k8[80]),
        .O(\a9/v1 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[16]_i_1__8 
       (.I0(k9[112]),
        .I1(k9[80]),
        .O(\a10/v1 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[17]_i_1 
       (.I0(k0[113]),
        .I1(k0[81]),
        .O(\a1/v1 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[17]_i_1__0 
       (.I0(k1[113]),
        .I1(k1[81]),
        .O(\a2/v1 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[17]_i_1__1 
       (.I0(k2[113]),
        .I1(k2[81]),
        .O(\a3/v1 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[17]_i_1__2 
       (.I0(k3[113]),
        .I1(k3[81]),
        .O(\a4/v1 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[17]_i_1__3 
       (.I0(k4[113]),
        .I1(k4[81]),
        .O(\a5/v1 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[17]_i_1__4 
       (.I0(k5[113]),
        .I1(k5[81]),
        .O(\a6/v1 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[17]_i_1__5 
       (.I0(k6[113]),
        .I1(k6[81]),
        .O(\a7/v1 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[17]_i_1__6 
       (.I0(k7[113]),
        .I1(k7[81]),
        .O(\a8/v1 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[17]_i_1__7 
       (.I0(k8[113]),
        .I1(k8[81]),
        .O(\a9/v1 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[17]_i_1__8 
       (.I0(k9[113]),
        .I1(k9[81]),
        .O(\a10/v1 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[18]_i_1 
       (.I0(k0[114]),
        .I1(k0[82]),
        .O(\a1/v1 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[18]_i_1__0 
       (.I0(k1[114]),
        .I1(k1[82]),
        .O(\a2/v1 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[18]_i_1__1 
       (.I0(k2[114]),
        .I1(k2[82]),
        .O(\a3/v1 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[18]_i_1__2 
       (.I0(k3[114]),
        .I1(k3[82]),
        .O(\a4/v1 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[18]_i_1__3 
       (.I0(k4[114]),
        .I1(k4[82]),
        .O(\a5/v1 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[18]_i_1__4 
       (.I0(k5[114]),
        .I1(k5[82]),
        .O(\a6/v1 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[18]_i_1__5 
       (.I0(k6[114]),
        .I1(k6[82]),
        .O(\a7/v1 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[18]_i_1__6 
       (.I0(k7[114]),
        .I1(k7[82]),
        .O(\a8/v1 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[18]_i_1__7 
       (.I0(k8[114]),
        .I1(k8[82]),
        .O(\a9/v1 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[18]_i_1__8 
       (.I0(k9[114]),
        .I1(k9[82]),
        .O(\a10/v1 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[19]_i_1 
       (.I0(k0[115]),
        .I1(k0[83]),
        .O(\a1/v1 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[19]_i_1__0 
       (.I0(k1[115]),
        .I1(k1[83]),
        .O(\a2/v1 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[19]_i_1__1 
       (.I0(k2[115]),
        .I1(k2[83]),
        .O(\a3/v1 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[19]_i_1__2 
       (.I0(k3[115]),
        .I1(k3[83]),
        .O(\a4/v1 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[19]_i_1__3 
       (.I0(k4[115]),
        .I1(k4[83]),
        .O(\a5/v1 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[19]_i_1__4 
       (.I0(k5[115]),
        .I1(k5[83]),
        .O(\a6/v1 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[19]_i_1__5 
       (.I0(k6[115]),
        .I1(k6[83]),
        .O(\a7/v1 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[19]_i_1__6 
       (.I0(k7[115]),
        .I1(k7[83]),
        .O(\a8/v1 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[19]_i_1__7 
       (.I0(k8[115]),
        .I1(k8[83]),
        .O(\a9/v1 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[19]_i_1__8 
       (.I0(k9[115]),
        .I1(k9[83]),
        .O(\a10/v1 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[1]_i_1 
       (.I0(k0[97]),
        .I1(k0[65]),
        .O(\a1/v1 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[1]_i_1__0 
       (.I0(k1[97]),
        .I1(k1[65]),
        .O(\a2/v1 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[1]_i_1__1 
       (.I0(k2[97]),
        .I1(k2[65]),
        .O(\a3/v1 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[1]_i_1__2 
       (.I0(k3[97]),
        .I1(k3[65]),
        .O(\a4/v1 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[1]_i_1__3 
       (.I0(k4[97]),
        .I1(k4[65]),
        .O(\a5/v1 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[1]_i_1__4 
       (.I0(k5[97]),
        .I1(k5[65]),
        .O(\a6/v1 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[1]_i_1__5 
       (.I0(k6[97]),
        .I1(k6[65]),
        .O(\a7/v1 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[1]_i_1__6 
       (.I0(k7[97]),
        .I1(k7[65]),
        .O(\a8/v1 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[1]_i_1__7 
       (.I0(k8[97]),
        .I1(k8[65]),
        .O(\a9/v1 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[1]_i_1__8 
       (.I0(k9[97]),
        .I1(k9[65]),
        .O(\a10/v1 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[20]_i_1 
       (.I0(k0[116]),
        .I1(k0[84]),
        .O(\a1/v1 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[20]_i_1__0 
       (.I0(k1[116]),
        .I1(k1[84]),
        .O(\a2/v1 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[20]_i_1__1 
       (.I0(k2[116]),
        .I1(k2[84]),
        .O(\a3/v1 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[20]_i_1__2 
       (.I0(k3[116]),
        .I1(k3[84]),
        .O(\a4/v1 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[20]_i_1__3 
       (.I0(k4[116]),
        .I1(k4[84]),
        .O(\a5/v1 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[20]_i_1__4 
       (.I0(k5[116]),
        .I1(k5[84]),
        .O(\a6/v1 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[20]_i_1__5 
       (.I0(k6[116]),
        .I1(k6[84]),
        .O(\a7/v1 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[20]_i_1__6 
       (.I0(k7[116]),
        .I1(k7[84]),
        .O(\a8/v1 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[20]_i_1__7 
       (.I0(k8[116]),
        .I1(k8[84]),
        .O(\a9/v1 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[20]_i_1__8 
       (.I0(k9[116]),
        .I1(k9[84]),
        .O(\a10/v1 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[21]_i_1 
       (.I0(k0[117]),
        .I1(k0[85]),
        .O(\a1/v1 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[21]_i_1__0 
       (.I0(k1[117]),
        .I1(k1[85]),
        .O(\a2/v1 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[21]_i_1__1 
       (.I0(k2[117]),
        .I1(k2[85]),
        .O(\a3/v1 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[21]_i_1__2 
       (.I0(k3[117]),
        .I1(k3[85]),
        .O(\a4/v1 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[21]_i_1__3 
       (.I0(k4[117]),
        .I1(k4[85]),
        .O(\a5/v1 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[21]_i_1__4 
       (.I0(k5[117]),
        .I1(k5[85]),
        .O(\a6/v1 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[21]_i_1__5 
       (.I0(k6[117]),
        .I1(k6[85]),
        .O(\a7/v1 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[21]_i_1__6 
       (.I0(k7[117]),
        .I1(k7[85]),
        .O(\a8/v1 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[21]_i_1__7 
       (.I0(k8[117]),
        .I1(k8[85]),
        .O(\a9/v1 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[21]_i_1__8 
       (.I0(k9[117]),
        .I1(k9[85]),
        .O(\a10/v1 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[22]_i_1 
       (.I0(k0[118]),
        .I1(k0[86]),
        .O(\a1/v1 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[22]_i_1__0 
       (.I0(k1[118]),
        .I1(k1[86]),
        .O(\a2/v1 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[22]_i_1__1 
       (.I0(k2[118]),
        .I1(k2[86]),
        .O(\a3/v1 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[22]_i_1__2 
       (.I0(k3[118]),
        .I1(k3[86]),
        .O(\a4/v1 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[22]_i_1__3 
       (.I0(k4[118]),
        .I1(k4[86]),
        .O(\a5/v1 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[22]_i_1__4 
       (.I0(k5[118]),
        .I1(k5[86]),
        .O(\a6/v1 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[22]_i_1__5 
       (.I0(k6[118]),
        .I1(k6[86]),
        .O(\a7/v1 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[22]_i_1__6 
       (.I0(k7[118]),
        .I1(k7[86]),
        .O(\a8/v1 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[22]_i_1__7 
       (.I0(k8[118]),
        .I1(k8[86]),
        .O(\a9/v1 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[22]_i_1__8 
       (.I0(k9[118]),
        .I1(k9[86]),
        .O(\a10/v1 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[23]_i_1 
       (.I0(k0[119]),
        .I1(k0[87]),
        .O(\a1/v1 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[23]_i_1__0 
       (.I0(k1[119]),
        .I1(k1[87]),
        .O(\a2/v1 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[23]_i_1__1 
       (.I0(k2[119]),
        .I1(k2[87]),
        .O(\a3/v1 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[23]_i_1__2 
       (.I0(k3[119]),
        .I1(k3[87]),
        .O(\a4/v1 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[23]_i_1__3 
       (.I0(k4[119]),
        .I1(k4[87]),
        .O(\a5/v1 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[23]_i_1__4 
       (.I0(k5[119]),
        .I1(k5[87]),
        .O(\a6/v1 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[23]_i_1__5 
       (.I0(k6[119]),
        .I1(k6[87]),
        .O(\a7/v1 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[23]_i_1__6 
       (.I0(k7[119]),
        .I1(k7[87]),
        .O(\a8/v1 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[23]_i_1__7 
       (.I0(k8[119]),
        .I1(k8[87]),
        .O(\a9/v1 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[23]_i_1__8 
       (.I0(k9[119]),
        .I1(k9[87]),
        .O(\a10/v1 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair879" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \k1a[24]_i_1 
       (.I0(k0[120]),
        .I1(k0[88]),
        .O(\k1a[24]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[24]_i_1__0 
       (.I0(k1[120]),
        .I1(k1[88]),
        .O(\a2/v1 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[24]_i_1__1 
       (.I0(k2[120]),
        .I1(k2[88]),
        .O(\a3/v1 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[24]_i_1__2 
       (.I0(k3[120]),
        .I1(k3[88]),
        .O(\a4/v1 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[24]_i_1__3 
       (.I0(k4[120]),
        .I1(k4[88]),
        .O(\a5/v1 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[24]_i_1__4 
       (.I0(k5[120]),
        .I1(k5[88]),
        .O(\a6/v1 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[24]_i_1__5 
       (.I0(k6[120]),
        .I1(k6[88]),
        .O(\a7/v1 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[24]_i_1__6 
       (.I0(k7[120]),
        .I1(k7[88]),
        .O(\a8/v1 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair451" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \k1a[24]_i_1__7 
       (.I0(k8[120]),
        .I1(k8[88]),
        .O(k1a));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[24]_i_1__8 
       (.I0(k9[120]),
        .I1(k9[88]),
        .O(\a10/v1 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[25]_i_1 
       (.I0(k0[121]),
        .I1(k0[89]),
        .O(\a1/v1 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair814" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \k1a[25]_i_1__0 
       (.I0(k1[121]),
        .I1(k1[89]),
        .O(\k1a[25]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[25]_i_1__1 
       (.I0(k2[121]),
        .I1(k2[89]),
        .O(\a3/v1 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[25]_i_1__2 
       (.I0(k3[121]),
        .I1(k3[89]),
        .O(\a4/v1 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[25]_i_1__3 
       (.I0(k4[121]),
        .I1(k4[89]),
        .O(\a5/v1 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[25]_i_1__4 
       (.I0(k5[121]),
        .I1(k5[89]),
        .O(\a6/v1 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[25]_i_1__5 
       (.I0(k6[121]),
        .I1(k6[89]),
        .O(\a7/v1 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[25]_i_1__6 
       (.I0(k7[121]),
        .I1(k7[89]),
        .O(\a8/v1 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair450" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \k1a[25]_i_1__7 
       (.I0(k8[121]),
        .I1(k8[89]),
        .O(\k1a[25]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair487" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \k1a[25]_i_1__8 
       (.I0(k9[121]),
        .I1(k9[89]),
        .O(\k1a[25]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[26]_i_1 
       (.I0(k0[122]),
        .I1(k0[90]),
        .O(\a1/v1 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[26]_i_1__0 
       (.I0(k1[122]),
        .I1(k1[90]),
        .O(\a2/v1 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair749" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \k1a[26]_i_1__1 
       (.I0(k2[122]),
        .I1(k2[90]),
        .O(\k1a[26]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[26]_i_1__2 
       (.I0(k3[122]),
        .I1(k3[90]),
        .O(\a4/v1 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[26]_i_1__3 
       (.I0(k4[122]),
        .I1(k4[90]),
        .O(\a5/v1 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[26]_i_1__4 
       (.I0(k5[122]),
        .I1(k5[90]),
        .O(\a6/v1 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[26]_i_1__5 
       (.I0(k6[122]),
        .I1(k6[90]),
        .O(\a7/v1 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[26]_i_1__6 
       (.I0(k7[122]),
        .I1(k7[90]),
        .O(\a8/v1 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[26]_i_1__7 
       (.I0(k8[122]),
        .I1(k8[90]),
        .O(\a9/v1 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair486" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \k1a[26]_i_1__8 
       (.I0(k9[122]),
        .I1(k9[90]),
        .O(\k1a[26]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[27]_i_1 
       (.I0(k0[123]),
        .I1(k0[91]),
        .O(\a1/v1 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[27]_i_1__0 
       (.I0(k1[123]),
        .I1(k1[91]),
        .O(\a2/v1 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[27]_i_1__1 
       (.I0(k2[123]),
        .I1(k2[91]),
        .O(\a3/v1 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair684" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \k1a[27]_i_1__2 
       (.I0(k3[123]),
        .I1(k3[91]),
        .O(\k1a[27]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[27]_i_1__3 
       (.I0(k4[123]),
        .I1(k4[91]),
        .O(\a5/v1 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[27]_i_1__4 
       (.I0(k5[123]),
        .I1(k5[91]),
        .O(\a6/v1 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[27]_i_1__5 
       (.I0(k6[123]),
        .I1(k6[91]),
        .O(\a7/v1 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[27]_i_1__6 
       (.I0(k7[123]),
        .I1(k7[91]),
        .O(\a8/v1 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair449" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \k1a[27]_i_1__7 
       (.I0(k8[123]),
        .I1(k8[91]),
        .O(\k1a[27]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[27]_i_1__8 
       (.I0(k9[123]),
        .I1(k9[91]),
        .O(\a10/v1 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[28]_i_1 
       (.I0(k0[124]),
        .I1(k0[92]),
        .O(\a1/v1 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[28]_i_1__0 
       (.I0(k1[124]),
        .I1(k1[92]),
        .O(\a2/v1 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[28]_i_1__1 
       (.I0(k2[124]),
        .I1(k2[92]),
        .O(\a3/v1 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[28]_i_1__2 
       (.I0(k3[124]),
        .I1(k3[92]),
        .O(\a4/v1 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair618" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \k1a[28]_i_1__3 
       (.I0(k4[124]),
        .I1(k4[92]),
        .O(\k1a[28]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[28]_i_1__4 
       (.I0(k5[124]),
        .I1(k5[92]),
        .O(\a6/v1 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[28]_i_1__5 
       (.I0(k6[124]),
        .I1(k6[92]),
        .O(\a7/v1 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[28]_i_1__6 
       (.I0(k7[124]),
        .I1(k7[92]),
        .O(\a8/v1 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair448" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \k1a[28]_i_1__7 
       (.I0(k8[124]),
        .I1(k8[92]),
        .O(\k1a[28]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair485" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \k1a[28]_i_1__8 
       (.I0(k9[124]),
        .I1(k9[92]),
        .O(\k1a[28]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[29]_i_1 
       (.I0(k0[125]),
        .I1(k0[93]),
        .O(\a1/v1 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[29]_i_1__0 
       (.I0(k1[125]),
        .I1(k1[93]),
        .O(\a2/v1 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[29]_i_1__1 
       (.I0(k2[125]),
        .I1(k2[93]),
        .O(\a3/v1 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[29]_i_1__2 
       (.I0(k3[125]),
        .I1(k3[93]),
        .O(\a4/v1 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[29]_i_1__3 
       (.I0(k4[125]),
        .I1(k4[93]),
        .O(\a5/v1 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair553" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \k1a[29]_i_1__4 
       (.I0(k5[125]),
        .I1(k5[93]),
        .O(\k1a[29]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[29]_i_1__5 
       (.I0(k6[125]),
        .I1(k6[93]),
        .O(\a7/v1 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[29]_i_1__6 
       (.I0(k7[125]),
        .I1(k7[93]),
        .O(\a8/v1 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[29]_i_1__7 
       (.I0(k8[125]),
        .I1(k8[93]),
        .O(\a9/v1 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair484" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \k1a[29]_i_1__8 
       (.I0(k9[125]),
        .I1(k9[93]),
        .O(\k1a[29]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[2]_i_1 
       (.I0(k0[98]),
        .I1(k0[66]),
        .O(\a1/v1 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[2]_i_1__0 
       (.I0(k1[98]),
        .I1(k1[66]),
        .O(\a2/v1 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[2]_i_1__1 
       (.I0(k2[98]),
        .I1(k2[66]),
        .O(\a3/v1 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[2]_i_1__2 
       (.I0(k3[98]),
        .I1(k3[66]),
        .O(\a4/v1 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[2]_i_1__3 
       (.I0(k4[98]),
        .I1(k4[66]),
        .O(\a5/v1 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[2]_i_1__4 
       (.I0(k5[98]),
        .I1(k5[66]),
        .O(\a6/v1 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[2]_i_1__5 
       (.I0(k6[98]),
        .I1(k6[66]),
        .O(\a7/v1 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[2]_i_1__6 
       (.I0(k7[98]),
        .I1(k7[66]),
        .O(\a8/v1 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[2]_i_1__7 
       (.I0(k8[98]),
        .I1(k8[66]),
        .O(\a9/v1 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[2]_i_1__8 
       (.I0(k9[98]),
        .I1(k9[66]),
        .O(\a10/v1 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[30]_i_1 
       (.I0(k0[126]),
        .I1(k0[94]),
        .O(\a1/v1 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[30]_i_1__0 
       (.I0(k1[126]),
        .I1(k1[94]),
        .O(\a2/v1 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[30]_i_1__1 
       (.I0(k2[126]),
        .I1(k2[94]),
        .O(\a3/v1 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[30]_i_1__2 
       (.I0(k3[126]),
        .I1(k3[94]),
        .O(\a4/v1 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[30]_i_1__3 
       (.I0(k4[126]),
        .I1(k4[94]),
        .O(\a5/v1 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[30]_i_1__4 
       (.I0(k5[126]),
        .I1(k5[94]),
        .O(\a6/v1 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair488" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \k1a[30]_i_1__5 
       (.I0(k6[126]),
        .I1(k6[94]),
        .O(\k1a[30]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[30]_i_1__6 
       (.I0(k7[126]),
        .I1(k7[94]),
        .O(\a8/v1 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[30]_i_1__7 
       (.I0(k8[126]),
        .I1(k8[94]),
        .O(\a9/v1 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[30]_i_1__8 
       (.I0(k9[126]),
        .I1(k9[94]),
        .O(\a10/v1 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[31]_i_1 
       (.I0(k0[127]),
        .I1(k0[95]),
        .O(\a1/v1 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[31]_i_1__0 
       (.I0(k1[127]),
        .I1(k1[95]),
        .O(\a2/v1 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[31]_i_1__1 
       (.I0(k2[127]),
        .I1(k2[95]),
        .O(\a3/v1 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[31]_i_1__2 
       (.I0(k3[127]),
        .I1(k3[95]),
        .O(\a4/v1 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[31]_i_1__3 
       (.I0(k4[127]),
        .I1(k4[95]),
        .O(\a5/v1 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[31]_i_1__4 
       (.I0(k5[127]),
        .I1(k5[95]),
        .O(\a6/v1 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[31]_i_1__5 
       (.I0(k6[127]),
        .I1(k6[95]),
        .O(\a7/v1 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair945" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \k1a[31]_i_1__6 
       (.I0(k7[127]),
        .I1(k7[95]),
        .O(\k1a[31]_i_1__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[31]_i_1__7 
       (.I0(k8[127]),
        .I1(k8[95]),
        .O(\a9/v1 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[31]_i_1__8 
       (.I0(k9[127]),
        .I1(k9[95]),
        .O(\a10/v1 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[3]_i_1 
       (.I0(k0[99]),
        .I1(k0[67]),
        .O(\a1/v1 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[3]_i_1__0 
       (.I0(k1[99]),
        .I1(k1[67]),
        .O(\a2/v1 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[3]_i_1__1 
       (.I0(k2[99]),
        .I1(k2[67]),
        .O(\a3/v1 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[3]_i_1__2 
       (.I0(k3[99]),
        .I1(k3[67]),
        .O(\a4/v1 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[3]_i_1__3 
       (.I0(k4[99]),
        .I1(k4[67]),
        .O(\a5/v1 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[3]_i_1__4 
       (.I0(k5[99]),
        .I1(k5[67]),
        .O(\a6/v1 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[3]_i_1__5 
       (.I0(k6[99]),
        .I1(k6[67]),
        .O(\a7/v1 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[3]_i_1__6 
       (.I0(k7[99]),
        .I1(k7[67]),
        .O(\a8/v1 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[3]_i_1__7 
       (.I0(k8[99]),
        .I1(k8[67]),
        .O(\a9/v1 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[3]_i_1__8 
       (.I0(k9[99]),
        .I1(k9[67]),
        .O(\a10/v1 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[4]_i_1 
       (.I0(k0[100]),
        .I1(k0[68]),
        .O(\a1/v1 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[4]_i_1__0 
       (.I0(k1[100]),
        .I1(k1[68]),
        .O(\a2/v1 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[4]_i_1__1 
       (.I0(k2[100]),
        .I1(k2[68]),
        .O(\a3/v1 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[4]_i_1__2 
       (.I0(k3[100]),
        .I1(k3[68]),
        .O(\a4/v1 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[4]_i_1__3 
       (.I0(k4[100]),
        .I1(k4[68]),
        .O(\a5/v1 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[4]_i_1__4 
       (.I0(k5[100]),
        .I1(k5[68]),
        .O(\a6/v1 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[4]_i_1__5 
       (.I0(k6[100]),
        .I1(k6[68]),
        .O(\a7/v1 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[4]_i_1__6 
       (.I0(k7[100]),
        .I1(k7[68]),
        .O(\a8/v1 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[4]_i_1__7 
       (.I0(k8[100]),
        .I1(k8[68]),
        .O(\a9/v1 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[4]_i_1__8 
       (.I0(k9[100]),
        .I1(k9[68]),
        .O(\a10/v1 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[5]_i_1 
       (.I0(k0[101]),
        .I1(k0[69]),
        .O(\a1/v1 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[5]_i_1__0 
       (.I0(k1[101]),
        .I1(k1[69]),
        .O(\a2/v1 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[5]_i_1__1 
       (.I0(k2[101]),
        .I1(k2[69]),
        .O(\a3/v1 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[5]_i_1__2 
       (.I0(k3[101]),
        .I1(k3[69]),
        .O(\a4/v1 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[5]_i_1__3 
       (.I0(k4[101]),
        .I1(k4[69]),
        .O(\a5/v1 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[5]_i_1__4 
       (.I0(k5[101]),
        .I1(k5[69]),
        .O(\a6/v1 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[5]_i_1__5 
       (.I0(k6[101]),
        .I1(k6[69]),
        .O(\a7/v1 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[5]_i_1__6 
       (.I0(k7[101]),
        .I1(k7[69]),
        .O(\a8/v1 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[5]_i_1__7 
       (.I0(k8[101]),
        .I1(k8[69]),
        .O(\a9/v1 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[5]_i_1__8 
       (.I0(k9[101]),
        .I1(k9[69]),
        .O(\a10/v1 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[6]_i_1 
       (.I0(k0[102]),
        .I1(k0[70]),
        .O(\a1/v1 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[6]_i_1__0 
       (.I0(k1[102]),
        .I1(k1[70]),
        .O(\a2/v1 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[6]_i_1__1 
       (.I0(k2[102]),
        .I1(k2[70]),
        .O(\a3/v1 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[6]_i_1__2 
       (.I0(k3[102]),
        .I1(k3[70]),
        .O(\a4/v1 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[6]_i_1__3 
       (.I0(k4[102]),
        .I1(k4[70]),
        .O(\a5/v1 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[6]_i_1__4 
       (.I0(k5[102]),
        .I1(k5[70]),
        .O(\a6/v1 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[6]_i_1__5 
       (.I0(k6[102]),
        .I1(k6[70]),
        .O(\a7/v1 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[6]_i_1__6 
       (.I0(k7[102]),
        .I1(k7[70]),
        .O(\a8/v1 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[6]_i_1__7 
       (.I0(k8[102]),
        .I1(k8[70]),
        .O(\a9/v1 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[6]_i_1__8 
       (.I0(k9[102]),
        .I1(k9[70]),
        .O(\a10/v1 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[7]_i_1 
       (.I0(k0[103]),
        .I1(k0[71]),
        .O(\a1/v1 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[7]_i_1__0 
       (.I0(k1[103]),
        .I1(k1[71]),
        .O(\a2/v1 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[7]_i_1__1 
       (.I0(k2[103]),
        .I1(k2[71]),
        .O(\a3/v1 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[7]_i_1__2 
       (.I0(k3[103]),
        .I1(k3[71]),
        .O(\a4/v1 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[7]_i_1__3 
       (.I0(k4[103]),
        .I1(k4[71]),
        .O(\a5/v1 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[7]_i_1__4 
       (.I0(k5[103]),
        .I1(k5[71]),
        .O(\a6/v1 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[7]_i_1__5 
       (.I0(k6[103]),
        .I1(k6[71]),
        .O(\a7/v1 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[7]_i_1__6 
       (.I0(k7[103]),
        .I1(k7[71]),
        .O(\a8/v1 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[7]_i_1__7 
       (.I0(k8[103]),
        .I1(k8[71]),
        .O(\a9/v1 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[7]_i_1__8 
       (.I0(k9[103]),
        .I1(k9[71]),
        .O(\a10/v1 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[8]_i_1 
       (.I0(k0[104]),
        .I1(k0[72]),
        .O(\a1/v1 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[8]_i_1__0 
       (.I0(k1[104]),
        .I1(k1[72]),
        .O(\a2/v1 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[8]_i_1__1 
       (.I0(k2[104]),
        .I1(k2[72]),
        .O(\a3/v1 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[8]_i_1__2 
       (.I0(k3[104]),
        .I1(k3[72]),
        .O(\a4/v1 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[8]_i_1__3 
       (.I0(k4[104]),
        .I1(k4[72]),
        .O(\a5/v1 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[8]_i_1__4 
       (.I0(k5[104]),
        .I1(k5[72]),
        .O(\a6/v1 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[8]_i_1__5 
       (.I0(k6[104]),
        .I1(k6[72]),
        .O(\a7/v1 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[8]_i_1__6 
       (.I0(k7[104]),
        .I1(k7[72]),
        .O(\a8/v1 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[8]_i_1__7 
       (.I0(k8[104]),
        .I1(k8[72]),
        .O(\a9/v1 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[8]_i_1__8 
       (.I0(k9[104]),
        .I1(k9[72]),
        .O(\a10/v1 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[9]_i_1 
       (.I0(k0[105]),
        .I1(k0[73]),
        .O(\a1/v1 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[9]_i_1__0 
       (.I0(k1[105]),
        .I1(k1[73]),
        .O(\a2/v1 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[9]_i_1__1 
       (.I0(k2[105]),
        .I1(k2[73]),
        .O(\a3/v1 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[9]_i_1__2 
       (.I0(k3[105]),
        .I1(k3[73]),
        .O(\a4/v1 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[9]_i_1__3 
       (.I0(k4[105]),
        .I1(k4[73]),
        .O(\a5/v1 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[9]_i_1__4 
       (.I0(k5[105]),
        .I1(k5[73]),
        .O(\a6/v1 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[9]_i_1__5 
       (.I0(k6[105]),
        .I1(k6[73]),
        .O(\a7/v1 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[9]_i_1__6 
       (.I0(k7[105]),
        .I1(k7[73]),
        .O(\a8/v1 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[9]_i_1__7 
       (.I0(k8[105]),
        .I1(k8[73]),
        .O(\a9/v1 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \k1a[9]_i_1__8 
       (.I0(k9[105]),
        .I1(k9[73]),
        .O(\a10/v1 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[0]_i_1 
       (.I0(k0[64]),
        .I1(k0[96]),
        .I2(k0[32]),
        .O(\a1/v2 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair101" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[0]_i_1__0 
       (.I0(k1[64]),
        .I1(k1[96]),
        .I2(k1[32]),
        .O(\a2/v2 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[0]_i_1__1 
       (.I0(k2[64]),
        .I1(k2[96]),
        .I2(k2[32]),
        .O(\a3/v2 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair26" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[0]_i_1__2 
       (.I0(k3[64]),
        .I1(k3[96]),
        .I2(k3[32]),
        .O(\a4/v2 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair9" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[0]_i_1__3 
       (.I0(k4[64]),
        .I1(k4[96]),
        .I2(k4[32]),
        .O(\a5/v2 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair36" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[0]_i_1__4 
       (.I0(k5[64]),
        .I1(k5[96]),
        .I2(k5[32]),
        .O(\a6/v2 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair261" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[0]_i_1__5 
       (.I0(k6[64]),
        .I1(k6[96]),
        .I2(k6[32]),
        .O(\a7/v2 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair316" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[0]_i_1__6 
       (.I0(k7[64]),
        .I1(k7[96]),
        .I2(k7[32]),
        .O(\a8/v2 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair192" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[0]_i_1__7 
       (.I0(k8[64]),
        .I1(k8[96]),
        .I2(k8[32]),
        .O(\a9/v2 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair223" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[0]_i_1__8 
       (.I0(k9[64]),
        .I1(k9[96]),
        .I2(k9[32]),
        .O(\a10/v2 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair183" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[10]_i_1 
       (.I0(k0[74]),
        .I1(k0[106]),
        .I2(k0[42]),
        .O(\a1/v2 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair154" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[10]_i_1__0 
       (.I0(k1[74]),
        .I1(k1[106]),
        .I2(k1[42]),
        .O(\a2/v2 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair125" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[10]_i_1__1 
       (.I0(k2[74]),
        .I1(k2[106]),
        .I2(k2[42]),
        .O(\a3/v2 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair92" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[10]_i_1__2 
       (.I0(k3[74]),
        .I1(k3[106]),
        .I2(k3[42]),
        .O(\a4/v2 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair33" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[10]_i_1__3 
       (.I0(k4[74]),
        .I1(k4[106]),
        .I2(k4[42]),
        .O(\a5/v2 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair46" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[10]_i_1__4 
       (.I0(k5[74]),
        .I1(k5[106]),
        .I2(k5[42]),
        .O(\a6/v2 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair271" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[10]_i_1__5 
       (.I0(k6[74]),
        .I1(k6[106]),
        .I2(k6[42]),
        .O(\a7/v2 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair306" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[10]_i_1__6 
       (.I0(k7[74]),
        .I1(k7[106]),
        .I2(k7[42]),
        .O(\a8/v2 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair201" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[10]_i_1__7 
       (.I0(k8[74]),
        .I1(k8[106]),
        .I2(k8[42]),
        .O(\a9/v2 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair233" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[10]_i_1__8 
       (.I0(k9[74]),
        .I1(k9[106]),
        .I2(k9[42]),
        .O(\a10/v2 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair182" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[11]_i_1 
       (.I0(k0[75]),
        .I1(k0[107]),
        .I2(k0[43]),
        .O(\a1/v2 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair153" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[11]_i_1__0 
       (.I0(k1[75]),
        .I1(k1[107]),
        .I2(k1[43]),
        .O(\a2/v2 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair124" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[11]_i_1__1 
       (.I0(k2[75]),
        .I1(k2[107]),
        .I2(k2[43]),
        .O(\a3/v2 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair91" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[11]_i_1__2 
       (.I0(k3[75]),
        .I1(k3[107]),
        .I2(k3[43]),
        .O(\a4/v2 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair32" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[11]_i_1__3 
       (.I0(k4[75]),
        .I1(k4[107]),
        .I2(k4[43]),
        .O(\a5/v2 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair47" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[11]_i_1__4 
       (.I0(k5[75]),
        .I1(k5[107]),
        .I2(k5[43]),
        .O(\a6/v2 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair272" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[11]_i_1__5 
       (.I0(k6[75]),
        .I1(k6[107]),
        .I2(k6[43]),
        .O(\a7/v2 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair305" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[11]_i_1__6 
       (.I0(k7[75]),
        .I1(k7[107]),
        .I2(k7[43]),
        .O(\a8/v2 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair202" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[11]_i_1__7 
       (.I0(k8[75]),
        .I1(k8[107]),
        .I2(k8[43]),
        .O(\a9/v2 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair234" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[11]_i_1__8 
       (.I0(k9[75]),
        .I1(k9[107]),
        .I2(k9[43]),
        .O(\a10/v2 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair181" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[12]_i_1 
       (.I0(k0[76]),
        .I1(k0[108]),
        .I2(k0[44]),
        .O(\a1/v2 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair152" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[12]_i_1__0 
       (.I0(k1[76]),
        .I1(k1[108]),
        .I2(k1[44]),
        .O(\a2/v2 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair123" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[12]_i_1__1 
       (.I0(k2[76]),
        .I1(k2[108]),
        .I2(k2[44]),
        .O(\a3/v2 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[12]_i_1__2 
       (.I0(k3[76]),
        .I1(k3[108]),
        .I2(k3[44]),
        .O(\a4/v2 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair31" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[12]_i_1__3 
       (.I0(k4[76]),
        .I1(k4[108]),
        .I2(k4[44]),
        .O(\a5/v2 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair48" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[12]_i_1__4 
       (.I0(k5[76]),
        .I1(k5[108]),
        .I2(k5[44]),
        .O(\a6/v2 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair273" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[12]_i_1__5 
       (.I0(k6[76]),
        .I1(k6[108]),
        .I2(k6[44]),
        .O(\a7/v2 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair304" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[12]_i_1__6 
       (.I0(k7[76]),
        .I1(k7[108]),
        .I2(k7[44]),
        .O(\a8/v2 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair203" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[12]_i_1__7 
       (.I0(k8[76]),
        .I1(k8[108]),
        .I2(k8[44]),
        .O(\a9/v2 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair235" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[12]_i_1__8 
       (.I0(k9[76]),
        .I1(k9[108]),
        .I2(k9[44]),
        .O(\a10/v2 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair180" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[13]_i_1 
       (.I0(k0[77]),
        .I1(k0[109]),
        .I2(k0[45]),
        .O(\a1/v2 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair151" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[13]_i_1__0 
       (.I0(k1[77]),
        .I1(k1[109]),
        .I2(k1[45]),
        .O(\a2/v2 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair122" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[13]_i_1__1 
       (.I0(k2[77]),
        .I1(k2[109]),
        .I2(k2[45]),
        .O(\a3/v2 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair89" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[13]_i_1__2 
       (.I0(k3[77]),
        .I1(k3[109]),
        .I2(k3[45]),
        .O(\a4/v2 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair30" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[13]_i_1__3 
       (.I0(k4[77]),
        .I1(k4[109]),
        .I2(k4[45]),
        .O(\a5/v2 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair49" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[13]_i_1__4 
       (.I0(k5[77]),
        .I1(k5[109]),
        .I2(k5[45]),
        .O(\a6/v2 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair274" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[13]_i_1__5 
       (.I0(k6[77]),
        .I1(k6[109]),
        .I2(k6[45]),
        .O(\a7/v2 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair303" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[13]_i_1__6 
       (.I0(k7[77]),
        .I1(k7[109]),
        .I2(k7[45]),
        .O(\a8/v2 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair204" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[13]_i_1__7 
       (.I0(k8[77]),
        .I1(k8[109]),
        .I2(k8[45]),
        .O(\a9/v2 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair236" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[13]_i_1__8 
       (.I0(k9[77]),
        .I1(k9[109]),
        .I2(k9[45]),
        .O(\a10/v2 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair179" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[14]_i_1 
       (.I0(k0[78]),
        .I1(k0[110]),
        .I2(k0[46]),
        .O(\a1/v2 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair150" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[14]_i_1__0 
       (.I0(k1[78]),
        .I1(k1[110]),
        .I2(k1[46]),
        .O(\a2/v2 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair121" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[14]_i_1__1 
       (.I0(k2[78]),
        .I1(k2[110]),
        .I2(k2[46]),
        .O(\a3/v2 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair88" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[14]_i_1__2 
       (.I0(k3[78]),
        .I1(k3[110]),
        .I2(k3[46]),
        .O(\a4/v2 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair29" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[14]_i_1__3 
       (.I0(k4[78]),
        .I1(k4[110]),
        .I2(k4[46]),
        .O(\a5/v2 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair50" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[14]_i_1__4 
       (.I0(k5[78]),
        .I1(k5[110]),
        .I2(k5[46]),
        .O(\a6/v2 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair275" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[14]_i_1__5 
       (.I0(k6[78]),
        .I1(k6[110]),
        .I2(k6[46]),
        .O(\a7/v2 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair302" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[14]_i_1__6 
       (.I0(k7[78]),
        .I1(k7[110]),
        .I2(k7[46]),
        .O(\a8/v2 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair205" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[14]_i_1__7 
       (.I0(k8[78]),
        .I1(k8[110]),
        .I2(k8[46]),
        .O(\a9/v2 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair237" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[14]_i_1__8 
       (.I0(k9[78]),
        .I1(k9[110]),
        .I2(k9[46]),
        .O(\a10/v2 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair178" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[15]_i_1 
       (.I0(k0[79]),
        .I1(k0[111]),
        .I2(k0[47]),
        .O(\a1/v2 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair149" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[15]_i_1__0 
       (.I0(k1[79]),
        .I1(k1[111]),
        .I2(k1[47]),
        .O(\a2/v2 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair120" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[15]_i_1__1 
       (.I0(k2[79]),
        .I1(k2[111]),
        .I2(k2[47]),
        .O(\a3/v2 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair87" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[15]_i_1__2 
       (.I0(k3[79]),
        .I1(k3[111]),
        .I2(k3[47]),
        .O(\a4/v2 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair28" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[15]_i_1__3 
       (.I0(k4[79]),
        .I1(k4[111]),
        .I2(k4[47]),
        .O(\a5/v2 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair51" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[15]_i_1__4 
       (.I0(k5[79]),
        .I1(k5[111]),
        .I2(k5[47]),
        .O(\a6/v2 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair276" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[15]_i_1__5 
       (.I0(k6[79]),
        .I1(k6[111]),
        .I2(k6[47]),
        .O(\a7/v2 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair301" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[15]_i_1__6 
       (.I0(k7[79]),
        .I1(k7[111]),
        .I2(k7[47]),
        .O(\a8/v2 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair206" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[15]_i_1__7 
       (.I0(k8[79]),
        .I1(k8[111]),
        .I2(k8[47]),
        .O(\a9/v2 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair238" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[15]_i_1__8 
       (.I0(k9[79]),
        .I1(k9[111]),
        .I2(k9[47]),
        .O(\a10/v2 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair177" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[16]_i_1 
       (.I0(k0[80]),
        .I1(k0[112]),
        .I2(k0[48]),
        .O(\a1/v2 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair148" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[16]_i_1__0 
       (.I0(k1[80]),
        .I1(k1[112]),
        .I2(k1[48]),
        .O(\a2/v2 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair119" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[16]_i_1__1 
       (.I0(k2[80]),
        .I1(k2[112]),
        .I2(k2[48]),
        .O(\a3/v2 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair86" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[16]_i_1__2 
       (.I0(k3[80]),
        .I1(k3[112]),
        .I2(k3[48]),
        .O(\a4/v2 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair27" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[16]_i_1__3 
       (.I0(k4[80]),
        .I1(k4[112]),
        .I2(k4[48]),
        .O(\a5/v2 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair52" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[16]_i_1__4 
       (.I0(k5[80]),
        .I1(k5[112]),
        .I2(k5[48]),
        .O(\a6/v2 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair277" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[16]_i_1__5 
       (.I0(k6[80]),
        .I1(k6[112]),
        .I2(k6[48]),
        .O(\a7/v2 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair300" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[16]_i_1__6 
       (.I0(k7[80]),
        .I1(k7[112]),
        .I2(k7[48]),
        .O(\a8/v2 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair207" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[16]_i_1__7 
       (.I0(k8[80]),
        .I1(k8[112]),
        .I2(k8[48]),
        .O(\a9/v2 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair239" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[16]_i_1__8 
       (.I0(k9[80]),
        .I1(k9[112]),
        .I2(k9[48]),
        .O(\a10/v2 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair176" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[17]_i_1 
       (.I0(k0[81]),
        .I1(k0[113]),
        .I2(k0[49]),
        .O(\a1/v2 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair147" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[17]_i_1__0 
       (.I0(k1[81]),
        .I1(k1[113]),
        .I2(k1[49]),
        .O(\a2/v2 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair118" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[17]_i_1__1 
       (.I0(k2[81]),
        .I1(k2[113]),
        .I2(k2[49]),
        .O(\a3/v2 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair85" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[17]_i_1__2 
       (.I0(k3[81]),
        .I1(k3[113]),
        .I2(k3[49]),
        .O(\a4/v2 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair102" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[17]_i_1__3 
       (.I0(k4[81]),
        .I1(k4[113]),
        .I2(k4[49]),
        .O(\a5/v2 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair53" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[17]_i_1__4 
       (.I0(k5[81]),
        .I1(k5[113]),
        .I2(k5[49]),
        .O(\a6/v2 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair278" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[17]_i_1__5 
       (.I0(k6[81]),
        .I1(k6[113]),
        .I2(k6[49]),
        .O(\a7/v2 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair299" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[17]_i_1__6 
       (.I0(k7[81]),
        .I1(k7[113]),
        .I2(k7[49]),
        .O(\a8/v2 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair208" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[17]_i_1__7 
       (.I0(k8[81]),
        .I1(k8[113]),
        .I2(k8[49]),
        .O(\a9/v2 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair240" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[17]_i_1__8 
       (.I0(k9[81]),
        .I1(k9[113]),
        .I2(k9[49]),
        .O(\a10/v2 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair175" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[18]_i_1 
       (.I0(k0[82]),
        .I1(k0[114]),
        .I2(k0[50]),
        .O(\a1/v2 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair146" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[18]_i_1__0 
       (.I0(k1[82]),
        .I1(k1[114]),
        .I2(k1[50]),
        .O(\a2/v2 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair117" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[18]_i_1__1 
       (.I0(k2[82]),
        .I1(k2[114]),
        .I2(k2[50]),
        .O(\a3/v2 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair84" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[18]_i_1__2 
       (.I0(k3[82]),
        .I1(k3[114]),
        .I2(k3[50]),
        .O(\a4/v2 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair25" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[18]_i_1__3 
       (.I0(k4[82]),
        .I1(k4[114]),
        .I2(k4[50]),
        .O(\a5/v2 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair54" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[18]_i_1__4 
       (.I0(k5[82]),
        .I1(k5[114]),
        .I2(k5[50]),
        .O(\a6/v2 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair279" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[18]_i_1__5 
       (.I0(k6[82]),
        .I1(k6[114]),
        .I2(k6[50]),
        .O(\a7/v2 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair298" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[18]_i_1__6 
       (.I0(k7[82]),
        .I1(k7[114]),
        .I2(k7[50]),
        .O(\a8/v2 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair209" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[18]_i_1__7 
       (.I0(k8[82]),
        .I1(k8[114]),
        .I2(k8[50]),
        .O(\a9/v2 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair241" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[18]_i_1__8 
       (.I0(k9[82]),
        .I1(k9[114]),
        .I2(k9[50]),
        .O(\a10/v2 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair174" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[19]_i_1 
       (.I0(k0[83]),
        .I1(k0[115]),
        .I2(k0[51]),
        .O(\a1/v2 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair145" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[19]_i_1__0 
       (.I0(k1[83]),
        .I1(k1[115]),
        .I2(k1[51]),
        .O(\a2/v2 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair116" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[19]_i_1__1 
       (.I0(k2[83]),
        .I1(k2[115]),
        .I2(k2[51]),
        .O(\a3/v2 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair83" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[19]_i_1__2 
       (.I0(k3[83]),
        .I1(k3[115]),
        .I2(k3[51]),
        .O(\a4/v2 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair24" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[19]_i_1__3 
       (.I0(k4[83]),
        .I1(k4[115]),
        .I2(k4[51]),
        .O(\a5/v2 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair55" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[19]_i_1__4 
       (.I0(k5[83]),
        .I1(k5[115]),
        .I2(k5[51]),
        .O(\a6/v2 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair280" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[19]_i_1__5 
       (.I0(k6[83]),
        .I1(k6[115]),
        .I2(k6[51]),
        .O(\a7/v2 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair297" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[19]_i_1__6 
       (.I0(k7[83]),
        .I1(k7[115]),
        .I2(k7[51]),
        .O(\a8/v2 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair210" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[19]_i_1__7 
       (.I0(k8[83]),
        .I1(k8[115]),
        .I2(k8[51]),
        .O(\a9/v2 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair242" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[19]_i_1__8 
       (.I0(k9[83]),
        .I1(k9[115]),
        .I2(k9[51]),
        .O(\a10/v2 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair103" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[1]_i_1 
       (.I0(k0[65]),
        .I1(k0[97]),
        .I2(k0[33]),
        .O(\a1/v2 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair11" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[1]_i_1__0 
       (.I0(k1[65]),
        .I1(k1[97]),
        .I2(k1[33]),
        .O(\a2/v2 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair10" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[1]_i_1__1 
       (.I0(k2[65]),
        .I1(k2[97]),
        .I2(k2[33]),
        .O(\a3/v2 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[1]_i_1__2 
       (.I0(k3[65]),
        .I1(k3[97]),
        .I2(k3[33]),
        .O(\a4/v2 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[1]_i_1__3 
       (.I0(k4[65]),
        .I1(k4[97]),
        .I2(k4[33]),
        .O(\a5/v2 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair37" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[1]_i_1__4 
       (.I0(k5[65]),
        .I1(k5[97]),
        .I2(k5[33]),
        .O(\a6/v2 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair262" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[1]_i_1__5 
       (.I0(k6[65]),
        .I1(k6[97]),
        .I2(k6[33]),
        .O(\a7/v2 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair315" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[1]_i_1__6 
       (.I0(k7[65]),
        .I1(k7[97]),
        .I2(k7[33]),
        .O(\a8/v2 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair318" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[1]_i_1__7 
       (.I0(k8[65]),
        .I1(k8[97]),
        .I2(k8[33]),
        .O(\a9/v2 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair224" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[1]_i_1__8 
       (.I0(k9[65]),
        .I1(k9[97]),
        .I2(k9[33]),
        .O(\a10/v2 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair173" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[20]_i_1 
       (.I0(k0[84]),
        .I1(k0[116]),
        .I2(k0[52]),
        .O(\a1/v2 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair144" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[20]_i_1__0 
       (.I0(k1[84]),
        .I1(k1[116]),
        .I2(k1[52]),
        .O(\a2/v2 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair115" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[20]_i_1__1 
       (.I0(k2[84]),
        .I1(k2[116]),
        .I2(k2[52]),
        .O(\a3/v2 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair82" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[20]_i_1__2 
       (.I0(k3[84]),
        .I1(k3[116]),
        .I2(k3[52]),
        .O(\a4/v2 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair23" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[20]_i_1__3 
       (.I0(k4[84]),
        .I1(k4[116]),
        .I2(k4[52]),
        .O(\a5/v2 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair56" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[20]_i_1__4 
       (.I0(k5[84]),
        .I1(k5[116]),
        .I2(k5[52]),
        .O(\a6/v2 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair281" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[20]_i_1__5 
       (.I0(k6[84]),
        .I1(k6[116]),
        .I2(k6[52]),
        .O(\a7/v2 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair296" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[20]_i_1__6 
       (.I0(k7[84]),
        .I1(k7[116]),
        .I2(k7[52]),
        .O(\a8/v2 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair211" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[20]_i_1__7 
       (.I0(k8[84]),
        .I1(k8[116]),
        .I2(k8[52]),
        .O(\a9/v2 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair243" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[20]_i_1__8 
       (.I0(k9[84]),
        .I1(k9[116]),
        .I2(k9[52]),
        .O(\a10/v2 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair172" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[21]_i_1 
       (.I0(k0[85]),
        .I1(k0[117]),
        .I2(k0[53]),
        .O(\a1/v2 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair143" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[21]_i_1__0 
       (.I0(k1[85]),
        .I1(k1[117]),
        .I2(k1[53]),
        .O(\a2/v2 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair114" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[21]_i_1__1 
       (.I0(k2[85]),
        .I1(k2[117]),
        .I2(k2[53]),
        .O(\a3/v2 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair81" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[21]_i_1__2 
       (.I0(k3[85]),
        .I1(k3[117]),
        .I2(k3[53]),
        .O(\a4/v2 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair22" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[21]_i_1__3 
       (.I0(k4[85]),
        .I1(k4[117]),
        .I2(k4[53]),
        .O(\a5/v2 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair57" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[21]_i_1__4 
       (.I0(k5[85]),
        .I1(k5[117]),
        .I2(k5[53]),
        .O(\a6/v2 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair282" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[21]_i_1__5 
       (.I0(k6[85]),
        .I1(k6[117]),
        .I2(k6[53]),
        .O(\a7/v2 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair295" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[21]_i_1__6 
       (.I0(k7[85]),
        .I1(k7[117]),
        .I2(k7[53]),
        .O(\a8/v2 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair212" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[21]_i_1__7 
       (.I0(k8[85]),
        .I1(k8[117]),
        .I2(k8[53]),
        .O(\a9/v2 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair244" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[21]_i_1__8 
       (.I0(k9[85]),
        .I1(k9[117]),
        .I2(k9[53]),
        .O(\a10/v2 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair171" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[22]_i_1 
       (.I0(k0[86]),
        .I1(k0[118]),
        .I2(k0[54]),
        .O(\a1/v2 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair142" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[22]_i_1__0 
       (.I0(k1[86]),
        .I1(k1[118]),
        .I2(k1[54]),
        .O(\a2/v2 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair113" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[22]_i_1__1 
       (.I0(k2[86]),
        .I1(k2[118]),
        .I2(k2[54]),
        .O(\a3/v2 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair80" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[22]_i_1__2 
       (.I0(k3[86]),
        .I1(k3[118]),
        .I2(k3[54]),
        .O(\a4/v2 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair21" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[22]_i_1__3 
       (.I0(k4[86]),
        .I1(k4[118]),
        .I2(k4[54]),
        .O(\a5/v2 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair58" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[22]_i_1__4 
       (.I0(k5[86]),
        .I1(k5[118]),
        .I2(k5[54]),
        .O(\a6/v2 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair283" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[22]_i_1__5 
       (.I0(k6[86]),
        .I1(k6[118]),
        .I2(k6[54]),
        .O(\a7/v2 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair294" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[22]_i_1__6 
       (.I0(k7[86]),
        .I1(k7[118]),
        .I2(k7[54]),
        .O(\a8/v2 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair213" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[22]_i_1__7 
       (.I0(k8[86]),
        .I1(k8[118]),
        .I2(k8[54]),
        .O(\a9/v2 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair245" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[22]_i_1__8 
       (.I0(k9[86]),
        .I1(k9[118]),
        .I2(k9[54]),
        .O(\a10/v2 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair170" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[23]_i_1 
       (.I0(k0[87]),
        .I1(k0[119]),
        .I2(k0[55]),
        .O(\a1/v2 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair141" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[23]_i_1__0 
       (.I0(k1[87]),
        .I1(k1[119]),
        .I2(k1[55]),
        .O(\a2/v2 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair112" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[23]_i_1__1 
       (.I0(k2[87]),
        .I1(k2[119]),
        .I2(k2[55]),
        .O(\a3/v2 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair79" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[23]_i_1__2 
       (.I0(k3[87]),
        .I1(k3[119]),
        .I2(k3[55]),
        .O(\a4/v2 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair20" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[23]_i_1__3 
       (.I0(k4[87]),
        .I1(k4[119]),
        .I2(k4[55]),
        .O(\a5/v2 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair59" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[23]_i_1__4 
       (.I0(k5[87]),
        .I1(k5[119]),
        .I2(k5[55]),
        .O(\a6/v2 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair284" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[23]_i_1__5 
       (.I0(k6[87]),
        .I1(k6[119]),
        .I2(k6[55]),
        .O(\a7/v2 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair317" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[23]_i_1__6 
       (.I0(k7[87]),
        .I1(k7[119]),
        .I2(k7[55]),
        .O(\a8/v2 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair214" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[23]_i_1__7 
       (.I0(k8[87]),
        .I1(k8[119]),
        .I2(k8[55]),
        .O(\a9/v2 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair246" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[23]_i_1__8 
       (.I0(k9[87]),
        .I1(k9[119]),
        .I2(k9[55]),
        .O(\a10/v2 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair162" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \k2a[24]_i_1 
       (.I0(k0[88]),
        .I1(k0[120]),
        .I2(k0[56]),
        .O(\a1/v2 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair140" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[24]_i_1__0 
       (.I0(k1[88]),
        .I1(k1[120]),
        .I2(k1[56]),
        .O(\a2/v2 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair111" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[24]_i_1__1 
       (.I0(k2[88]),
        .I1(k2[120]),
        .I2(k2[56]),
        .O(\a3/v2 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair78" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[24]_i_1__2 
       (.I0(k3[88]),
        .I1(k3[120]),
        .I2(k3[56]),
        .O(\a4/v2 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair19" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[24]_i_1__3 
       (.I0(k4[88]),
        .I1(k4[120]),
        .I2(k4[56]),
        .O(\a5/v2 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair60" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[24]_i_1__4 
       (.I0(k5[88]),
        .I1(k5[120]),
        .I2(k5[56]),
        .O(\a6/v2 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair285" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[24]_i_1__5 
       (.I0(k6[88]),
        .I1(k6[120]),
        .I2(k6[56]),
        .O(\a7/v2 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair260" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[24]_i_1__6 
       (.I0(k7[88]),
        .I1(k7[120]),
        .I2(k7[56]),
        .O(\a8/v2 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair219" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \k2a[24]_i_1__7 
       (.I0(k8[88]),
        .I1(k8[120]),
        .I2(k8[56]),
        .O(\a9/v2 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair247" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[24]_i_1__8 
       (.I0(k9[88]),
        .I1(k9[120]),
        .I2(k9[56]),
        .O(\a10/v2 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair169" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[25]_i_1 
       (.I0(k0[89]),
        .I1(k0[121]),
        .I2(k0[57]),
        .O(\a1/v2 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair133" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \k2a[25]_i_1__0 
       (.I0(k1[89]),
        .I1(k1[121]),
        .I2(k1[57]),
        .O(\a2/v2 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair110" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[25]_i_1__1 
       (.I0(k2[89]),
        .I1(k2[121]),
        .I2(k2[57]),
        .O(\a3/v2 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair77" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[25]_i_1__2 
       (.I0(k3[89]),
        .I1(k3[121]),
        .I2(k3[57]),
        .O(\a4/v2 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair18" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[25]_i_1__3 
       (.I0(k4[89]),
        .I1(k4[121]),
        .I2(k4[57]),
        .O(\a5/v2 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair61" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[25]_i_1__4 
       (.I0(k5[89]),
        .I1(k5[121]),
        .I2(k5[57]),
        .O(\a6/v2 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair286" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[25]_i_1__5 
       (.I0(k6[89]),
        .I1(k6[121]),
        .I2(k6[57]),
        .O(\a7/v2 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair259" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[25]_i_1__6 
       (.I0(k7[89]),
        .I1(k7[121]),
        .I2(k7[57]),
        .O(\a8/v2 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair220" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \k2a[25]_i_1__7 
       (.I0(k8[89]),
        .I1(k8[121]),
        .I2(k8[57]),
        .O(\a9/v2 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair251" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \k2a[25]_i_1__8 
       (.I0(k9[89]),
        .I1(k9[121]),
        .I2(k9[57]),
        .O(\a10/v2 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair168" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[26]_i_1 
       (.I0(k0[90]),
        .I1(k0[122]),
        .I2(k0[58]),
        .O(\a1/v2 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair139" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[26]_i_1__0 
       (.I0(k1[90]),
        .I1(k1[122]),
        .I2(k1[58]),
        .O(\a2/v2 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair104" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \k2a[26]_i_1__1 
       (.I0(k2[90]),
        .I1(k2[122]),
        .I2(k2[58]),
        .O(\a3/v2 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair76" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[26]_i_1__2 
       (.I0(k3[90]),
        .I1(k3[122]),
        .I2(k3[58]),
        .O(\a4/v2 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair17" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[26]_i_1__3 
       (.I0(k4[90]),
        .I1(k4[122]),
        .I2(k4[58]),
        .O(\a5/v2 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair62" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[26]_i_1__4 
       (.I0(k5[90]),
        .I1(k5[122]),
        .I2(k5[58]),
        .O(\a6/v2 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair287" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[26]_i_1__5 
       (.I0(k6[90]),
        .I1(k6[122]),
        .I2(k6[58]),
        .O(\a7/v2 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair258" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[26]_i_1__6 
       (.I0(k7[90]),
        .I1(k7[122]),
        .I2(k7[58]),
        .O(\a8/v2 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair215" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[26]_i_1__7 
       (.I0(k8[90]),
        .I1(k8[122]),
        .I2(k8[58]),
        .O(\a9/v2 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair252" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \k2a[26]_i_1__8 
       (.I0(k9[90]),
        .I1(k9[122]),
        .I2(k9[58]),
        .O(\a10/v2 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair167" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[27]_i_1 
       (.I0(k0[91]),
        .I1(k0[123]),
        .I2(k0[59]),
        .O(\a1/v2 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair138" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[27]_i_1__0 
       (.I0(k1[91]),
        .I1(k1[123]),
        .I2(k1[59]),
        .O(\a2/v2 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair109" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[27]_i_1__1 
       (.I0(k2[91]),
        .I1(k2[123]),
        .I2(k2[59]),
        .O(\a3/v2 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair71" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \k2a[27]_i_1__2 
       (.I0(k3[91]),
        .I1(k3[123]),
        .I2(k3[59]),
        .O(\a4/v2 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair16" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[27]_i_1__3 
       (.I0(k4[91]),
        .I1(k4[123]),
        .I2(k4[59]),
        .O(\a5/v2 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair63" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[27]_i_1__4 
       (.I0(k5[91]),
        .I1(k5[123]),
        .I2(k5[59]),
        .O(\a6/v2 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair288" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[27]_i_1__5 
       (.I0(k6[91]),
        .I1(k6[123]),
        .I2(k6[59]),
        .O(\a7/v2 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair257" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[27]_i_1__6 
       (.I0(k7[91]),
        .I1(k7[123]),
        .I2(k7[59]),
        .O(\a8/v2 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair221" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \k2a[27]_i_1__7 
       (.I0(k8[91]),
        .I1(k8[123]),
        .I2(k8[59]),
        .O(\a9/v2 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair248" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[27]_i_1__8 
       (.I0(k9[91]),
        .I1(k9[123]),
        .I2(k9[59]),
        .O(\a10/v2 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair166" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[28]_i_1 
       (.I0(k0[92]),
        .I1(k0[124]),
        .I2(k0[60]),
        .O(\a1/v2 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair137" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[28]_i_1__0 
       (.I0(k1[92]),
        .I1(k1[124]),
        .I2(k1[60]),
        .O(\a2/v2 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair108" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[28]_i_1__1 
       (.I0(k2[92]),
        .I1(k2[124]),
        .I2(k2[60]),
        .O(\a3/v2 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair75" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[28]_i_1__2 
       (.I0(k3[92]),
        .I1(k3[124]),
        .I2(k3[60]),
        .O(\a4/v2 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair12" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \k2a[28]_i_1__3 
       (.I0(k4[92]),
        .I1(k4[124]),
        .I2(k4[60]),
        .O(\a5/v2 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair64" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[28]_i_1__4 
       (.I0(k5[92]),
        .I1(k5[124]),
        .I2(k5[60]),
        .O(\a6/v2 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair289" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[28]_i_1__5 
       (.I0(k6[92]),
        .I1(k6[124]),
        .I2(k6[60]),
        .O(\a7/v2 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair256" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[28]_i_1__6 
       (.I0(k7[92]),
        .I1(k7[124]),
        .I2(k7[60]),
        .O(\a8/v2 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair222" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \k2a[28]_i_1__7 
       (.I0(k8[92]),
        .I1(k8[124]),
        .I2(k8[60]),
        .O(\a9/v2 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair253" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \k2a[28]_i_1__8 
       (.I0(k9[92]),
        .I1(k9[124]),
        .I2(k9[60]),
        .O(\a10/v2 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair165" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[29]_i_1 
       (.I0(k0[93]),
        .I1(k0[125]),
        .I2(k0[61]),
        .O(\a1/v2 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair136" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[29]_i_1__0 
       (.I0(k1[93]),
        .I1(k1[125]),
        .I2(k1[61]),
        .O(\a2/v2 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair107" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[29]_i_1__1 
       (.I0(k2[93]),
        .I1(k2[125]),
        .I2(k2[61]),
        .O(\a3/v2 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair74" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[29]_i_1__2 
       (.I0(k3[93]),
        .I1(k3[125]),
        .I2(k3[61]),
        .O(\a4/v2 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair15" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[29]_i_1__3 
       (.I0(k4[93]),
        .I1(k4[125]),
        .I2(k4[61]),
        .O(\a5/v2 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair67" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \k2a[29]_i_1__4 
       (.I0(k5[93]),
        .I1(k5[125]),
        .I2(k5[61]),
        .O(\a6/v2 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair290" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[29]_i_1__5 
       (.I0(k6[93]),
        .I1(k6[125]),
        .I2(k6[61]),
        .O(\a7/v2 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair255" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[29]_i_1__6 
       (.I0(k7[93]),
        .I1(k7[125]),
        .I2(k7[61]),
        .O(\a8/v2 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair216" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[29]_i_1__7 
       (.I0(k8[93]),
        .I1(k8[125]),
        .I2(k8[61]),
        .O(\a9/v2 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair254" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \k2a[29]_i_1__8 
       (.I0(k9[93]),
        .I1(k9[125]),
        .I2(k9[61]),
        .O(\a10/v2 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair191" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[2]_i_1 
       (.I0(k0[66]),
        .I1(k0[98]),
        .I2(k0[34]),
        .O(\a1/v2 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[2]_i_1__0 
       (.I0(k1[66]),
        .I1(k1[98]),
        .I2(k1[34]),
        .O(\a2/v2 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[2]_i_1__1 
       (.I0(k2[66]),
        .I1(k2[98]),
        .I2(k2[34]),
        .O(\a3/v2 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair100" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[2]_i_1__2 
       (.I0(k3[66]),
        .I1(k3[98]),
        .I2(k3[34]),
        .O(\a4/v2 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair35" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[2]_i_1__3 
       (.I0(k4[66]),
        .I1(k4[98]),
        .I2(k4[34]),
        .O(\a5/v2 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair38" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[2]_i_1__4 
       (.I0(k5[66]),
        .I1(k5[98]),
        .I2(k5[34]),
        .O(\a6/v2 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair263" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[2]_i_1__5 
       (.I0(k6[66]),
        .I1(k6[98]),
        .I2(k6[34]),
        .O(\a7/v2 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair314" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[2]_i_1__6 
       (.I0(k7[66]),
        .I1(k7[98]),
        .I2(k7[34]),
        .O(\a8/v2 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair193" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[2]_i_1__7 
       (.I0(k8[66]),
        .I1(k8[98]),
        .I2(k8[34]),
        .O(\a9/v2 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair225" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[2]_i_1__8 
       (.I0(k9[66]),
        .I1(k9[98]),
        .I2(k9[34]),
        .O(\a10/v2 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair164" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[30]_i_1 
       (.I0(k0[94]),
        .I1(k0[126]),
        .I2(k0[62]),
        .O(\a1/v2 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair135" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[30]_i_1__0 
       (.I0(k1[94]),
        .I1(k1[126]),
        .I2(k1[62]),
        .O(\a2/v2 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair106" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[30]_i_1__1 
       (.I0(k2[94]),
        .I1(k2[126]),
        .I2(k2[62]),
        .O(\a3/v2 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair73" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[30]_i_1__2 
       (.I0(k3[94]),
        .I1(k3[126]),
        .I2(k3[62]),
        .O(\a4/v2 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[30]_i_1__3 
       (.I0(k4[94]),
        .I1(k4[126]),
        .I2(k4[62]),
        .O(\a5/v2 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair65" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[30]_i_1__4 
       (.I0(k5[94]),
        .I1(k5[126]),
        .I2(k5[62]),
        .O(\a6/v2 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair292" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \k2a[30]_i_1__5 
       (.I0(k6[94]),
        .I1(k6[126]),
        .I2(k6[62]),
        .O(\a7/v2 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair293" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[30]_i_1__6 
       (.I0(k7[94]),
        .I1(k7[126]),
        .I2(k7[62]),
        .O(\a8/v2 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair217" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[30]_i_1__7 
       (.I0(k8[94]),
        .I1(k8[126]),
        .I2(k8[62]),
        .O(\a9/v2 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair249" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[30]_i_1__8 
       (.I0(k9[94]),
        .I1(k9[126]),
        .I2(k9[62]),
        .O(\a10/v2 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair163" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[31]_i_1 
       (.I0(k0[95]),
        .I1(k0[127]),
        .I2(k0[63]),
        .O(\a1/v2 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair134" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[31]_i_1__0 
       (.I0(k1[95]),
        .I1(k1[127]),
        .I2(k1[63]),
        .O(\a2/v2 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair105" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[31]_i_1__1 
       (.I0(k2[95]),
        .I1(k2[127]),
        .I2(k2[63]),
        .O(\a3/v2 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair72" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[31]_i_1__2 
       (.I0(k3[95]),
        .I1(k3[127]),
        .I2(k3[63]),
        .O(\a4/v2 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[31]_i_1__3 
       (.I0(k4[95]),
        .I1(k4[127]),
        .I2(k4[63]),
        .O(\a5/v2 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair66" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[31]_i_1__4 
       (.I0(k5[95]),
        .I1(k5[127]),
        .I2(k5[63]),
        .O(\a6/v2 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair291" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[31]_i_1__5 
       (.I0(k6[95]),
        .I1(k6[127]),
        .I2(k6[63]),
        .O(\a7/v2 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair319" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \k2a[31]_i_1__6 
       (.I0(k7[95]),
        .I1(k7[127]),
        .I2(k7[63]),
        .O(\a8/v2 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair218" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[31]_i_1__7 
       (.I0(k8[95]),
        .I1(k8[127]),
        .I2(k8[63]),
        .O(\a9/v2 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair250" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[31]_i_1__8 
       (.I0(k9[95]),
        .I1(k9[127]),
        .I2(k9[63]),
        .O(\a10/v2 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair190" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[3]_i_1 
       (.I0(k0[67]),
        .I1(k0[99]),
        .I2(k0[35]),
        .O(\a1/v2 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair161" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[3]_i_1__0 
       (.I0(k1[67]),
        .I1(k1[99]),
        .I2(k1[35]),
        .O(\a2/v2 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair132" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[3]_i_1__1 
       (.I0(k2[67]),
        .I1(k2[99]),
        .I2(k2[35]),
        .O(\a3/v2 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair99" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[3]_i_1__2 
       (.I0(k3[67]),
        .I1(k3[99]),
        .I2(k3[35]),
        .O(\a4/v2 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair70" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[3]_i_1__3 
       (.I0(k4[67]),
        .I1(k4[99]),
        .I2(k4[35]),
        .O(\a5/v2 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair39" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[3]_i_1__4 
       (.I0(k5[67]),
        .I1(k5[99]),
        .I2(k5[35]),
        .O(\a6/v2 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair264" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[3]_i_1__5 
       (.I0(k6[67]),
        .I1(k6[99]),
        .I2(k6[35]),
        .O(\a7/v2 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair313" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[3]_i_1__6 
       (.I0(k7[67]),
        .I1(k7[99]),
        .I2(k7[35]),
        .O(\a8/v2 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair194" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[3]_i_1__7 
       (.I0(k8[67]),
        .I1(k8[99]),
        .I2(k8[35]),
        .O(\a9/v2 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair226" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[3]_i_1__8 
       (.I0(k9[67]),
        .I1(k9[99]),
        .I2(k9[35]),
        .O(\a10/v2 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair189" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[4]_i_1 
       (.I0(k0[68]),
        .I1(k0[100]),
        .I2(k0[36]),
        .O(\a1/v2 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair160" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[4]_i_1__0 
       (.I0(k1[68]),
        .I1(k1[100]),
        .I2(k1[36]),
        .O(\a2/v2 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair131" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[4]_i_1__1 
       (.I0(k2[68]),
        .I1(k2[100]),
        .I2(k2[36]),
        .O(\a3/v2 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair98" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[4]_i_1__2 
       (.I0(k3[68]),
        .I1(k3[100]),
        .I2(k3[36]),
        .O(\a4/v2 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair69" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[4]_i_1__3 
       (.I0(k4[68]),
        .I1(k4[100]),
        .I2(k4[36]),
        .O(\a5/v2 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair40" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[4]_i_1__4 
       (.I0(k5[68]),
        .I1(k5[100]),
        .I2(k5[36]),
        .O(\a6/v2 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair265" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[4]_i_1__5 
       (.I0(k6[68]),
        .I1(k6[100]),
        .I2(k6[36]),
        .O(\a7/v2 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair312" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[4]_i_1__6 
       (.I0(k7[68]),
        .I1(k7[100]),
        .I2(k7[36]),
        .O(\a8/v2 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair195" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[4]_i_1__7 
       (.I0(k8[68]),
        .I1(k8[100]),
        .I2(k8[36]),
        .O(\a9/v2 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair227" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[4]_i_1__8 
       (.I0(k9[68]),
        .I1(k9[100]),
        .I2(k9[36]),
        .O(\a10/v2 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair188" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[5]_i_1 
       (.I0(k0[69]),
        .I1(k0[101]),
        .I2(k0[37]),
        .O(\a1/v2 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair159" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[5]_i_1__0 
       (.I0(k1[69]),
        .I1(k1[101]),
        .I2(k1[37]),
        .O(\a2/v2 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair130" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[5]_i_1__1 
       (.I0(k2[69]),
        .I1(k2[101]),
        .I2(k2[37]),
        .O(\a3/v2 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair97" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[5]_i_1__2 
       (.I0(k3[69]),
        .I1(k3[101]),
        .I2(k3[37]),
        .O(\a4/v2 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair68" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[5]_i_1__3 
       (.I0(k4[69]),
        .I1(k4[101]),
        .I2(k4[37]),
        .O(\a5/v2 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair41" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[5]_i_1__4 
       (.I0(k5[69]),
        .I1(k5[101]),
        .I2(k5[37]),
        .O(\a6/v2 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair266" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[5]_i_1__5 
       (.I0(k6[69]),
        .I1(k6[101]),
        .I2(k6[37]),
        .O(\a7/v2 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair311" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[5]_i_1__6 
       (.I0(k7[69]),
        .I1(k7[101]),
        .I2(k7[37]),
        .O(\a8/v2 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair196" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[5]_i_1__7 
       (.I0(k8[69]),
        .I1(k8[101]),
        .I2(k8[37]),
        .O(\a9/v2 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair228" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[5]_i_1__8 
       (.I0(k9[69]),
        .I1(k9[101]),
        .I2(k9[37]),
        .O(\a10/v2 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair187" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[6]_i_1 
       (.I0(k0[70]),
        .I1(k0[102]),
        .I2(k0[38]),
        .O(\a1/v2 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair158" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[6]_i_1__0 
       (.I0(k1[70]),
        .I1(k1[102]),
        .I2(k1[38]),
        .O(\a2/v2 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair129" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[6]_i_1__1 
       (.I0(k2[70]),
        .I1(k2[102]),
        .I2(k2[38]),
        .O(\a3/v2 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair96" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[6]_i_1__2 
       (.I0(k3[70]),
        .I1(k3[102]),
        .I2(k3[38]),
        .O(\a4/v2 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[6]_i_1__3 
       (.I0(k4[70]),
        .I1(k4[102]),
        .I2(k4[38]),
        .O(\a5/v2 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair42" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[6]_i_1__4 
       (.I0(k5[70]),
        .I1(k5[102]),
        .I2(k5[38]),
        .O(\a6/v2 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair267" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[6]_i_1__5 
       (.I0(k6[70]),
        .I1(k6[102]),
        .I2(k6[38]),
        .O(\a7/v2 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair310" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[6]_i_1__6 
       (.I0(k7[70]),
        .I1(k7[102]),
        .I2(k7[38]),
        .O(\a8/v2 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair197" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[6]_i_1__7 
       (.I0(k8[70]),
        .I1(k8[102]),
        .I2(k8[38]),
        .O(\a9/v2 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair229" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[6]_i_1__8 
       (.I0(k9[70]),
        .I1(k9[102]),
        .I2(k9[38]),
        .O(\a10/v2 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair186" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[7]_i_1 
       (.I0(k0[71]),
        .I1(k0[103]),
        .I2(k0[39]),
        .O(\a1/v2 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair157" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[7]_i_1__0 
       (.I0(k1[71]),
        .I1(k1[103]),
        .I2(k1[39]),
        .O(\a2/v2 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair128" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[7]_i_1__1 
       (.I0(k2[71]),
        .I1(k2[103]),
        .I2(k2[39]),
        .O(\a3/v2 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair95" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[7]_i_1__2 
       (.I0(k3[71]),
        .I1(k3[103]),
        .I2(k3[39]),
        .O(\a4/v2 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair1" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[7]_i_1__3 
       (.I0(k4[71]),
        .I1(k4[103]),
        .I2(k4[39]),
        .O(\a5/v2 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair43" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[7]_i_1__4 
       (.I0(k5[71]),
        .I1(k5[103]),
        .I2(k5[39]),
        .O(\a6/v2 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair268" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[7]_i_1__5 
       (.I0(k6[71]),
        .I1(k6[103]),
        .I2(k6[39]),
        .O(\a7/v2 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair309" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[7]_i_1__6 
       (.I0(k7[71]),
        .I1(k7[103]),
        .I2(k7[39]),
        .O(\a8/v2 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair198" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[7]_i_1__7 
       (.I0(k8[71]),
        .I1(k8[103]),
        .I2(k8[39]),
        .O(\a9/v2 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair230" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[7]_i_1__8 
       (.I0(k9[71]),
        .I1(k9[103]),
        .I2(k9[39]),
        .O(\a10/v2 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair185" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[8]_i_1 
       (.I0(k0[72]),
        .I1(k0[104]),
        .I2(k0[40]),
        .O(\a1/v2 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair156" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[8]_i_1__0 
       (.I0(k1[72]),
        .I1(k1[104]),
        .I2(k1[40]),
        .O(\a2/v2 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair127" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[8]_i_1__1 
       (.I0(k2[72]),
        .I1(k2[104]),
        .I2(k2[40]),
        .O(\a3/v2 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair94" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[8]_i_1__2 
       (.I0(k3[72]),
        .I1(k3[104]),
        .I2(k3[40]),
        .O(\a4/v2 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair0" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[8]_i_1__3 
       (.I0(k4[72]),
        .I1(k4[104]),
        .I2(k4[40]),
        .O(\a5/v2 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair44" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[8]_i_1__4 
       (.I0(k5[72]),
        .I1(k5[104]),
        .I2(k5[40]),
        .O(\a6/v2 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair269" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[8]_i_1__5 
       (.I0(k6[72]),
        .I1(k6[104]),
        .I2(k6[40]),
        .O(\a7/v2 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair308" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[8]_i_1__6 
       (.I0(k7[72]),
        .I1(k7[104]),
        .I2(k7[40]),
        .O(\a8/v2 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair199" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[8]_i_1__7 
       (.I0(k8[72]),
        .I1(k8[104]),
        .I2(k8[40]),
        .O(\a9/v2 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair231" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[8]_i_1__8 
       (.I0(k9[72]),
        .I1(k9[104]),
        .I2(k9[40]),
        .O(\a10/v2 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair184" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[9]_i_1 
       (.I0(k0[73]),
        .I1(k0[105]),
        .I2(k0[41]),
        .O(\a1/v2 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair155" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[9]_i_1__0 
       (.I0(k1[73]),
        .I1(k1[105]),
        .I2(k1[41]),
        .O(\a2/v2 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair126" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[9]_i_1__1 
       (.I0(k2[73]),
        .I1(k2[105]),
        .I2(k2[41]),
        .O(\a3/v2 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair93" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[9]_i_1__2 
       (.I0(k3[73]),
        .I1(k3[105]),
        .I2(k3[41]),
        .O(\a4/v2 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair34" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[9]_i_1__3 
       (.I0(k4[73]),
        .I1(k4[105]),
        .I2(k4[41]),
        .O(\a5/v2 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair45" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[9]_i_1__4 
       (.I0(k5[73]),
        .I1(k5[105]),
        .I2(k5[41]),
        .O(\a6/v2 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair270" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[9]_i_1__5 
       (.I0(k6[73]),
        .I1(k6[105]),
        .I2(k6[41]),
        .O(\a7/v2 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair307" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[9]_i_1__6 
       (.I0(k7[73]),
        .I1(k7[105]),
        .I2(k7[41]),
        .O(\a8/v2 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair200" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[9]_i_1__7 
       (.I0(k8[73]),
        .I1(k8[105]),
        .I2(k8[41]),
        .O(\a9/v2 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair232" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \k2a[9]_i_1__8 
       (.I0(k9[73]),
        .I1(k9[105]),
        .I2(k9[41]),
        .O(\a10/v2 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[0]_i_1 
       (.I0(k0[32]),
        .I1(k0[96]),
        .I2(k0[64]),
        .I3(k0[0]),
        .O(\a1/v3 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair101" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[0]_i_1__0 
       (.I0(k1[32]),
        .I1(k1[96]),
        .I2(k1[64]),
        .I3(k1[0]),
        .O(\a2/v3 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[0]_i_1__1 
       (.I0(k2[32]),
        .I1(k2[96]),
        .I2(k2[64]),
        .I3(k2[0]),
        .O(\a3/v3 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair26" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[0]_i_1__2 
       (.I0(k3[32]),
        .I1(k3[96]),
        .I2(k3[64]),
        .I3(k3[0]),
        .O(\a4/v3 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair9" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[0]_i_1__3 
       (.I0(k4[32]),
        .I1(k4[96]),
        .I2(k4[64]),
        .I3(k4[0]),
        .O(\a5/v3 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair36" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[0]_i_1__4 
       (.I0(k5[32]),
        .I1(k5[96]),
        .I2(k5[64]),
        .I3(k5[0]),
        .O(\a6/v3 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair261" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[0]_i_1__5 
       (.I0(k6[32]),
        .I1(k6[96]),
        .I2(k6[64]),
        .I3(k6[0]),
        .O(\a7/v3 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair316" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[0]_i_1__6 
       (.I0(k7[32]),
        .I1(k7[96]),
        .I2(k7[64]),
        .I3(k7[0]),
        .O(\a8/v3 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair192" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[0]_i_1__7 
       (.I0(k8[32]),
        .I1(k8[96]),
        .I2(k8[64]),
        .I3(k8[0]),
        .O(\a9/v3 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair223" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[0]_i_1__8 
       (.I0(k9[32]),
        .I1(k9[96]),
        .I2(k9[64]),
        .I3(k9[0]),
        .O(\a10/v3 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair183" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[10]_i_1 
       (.I0(k0[42]),
        .I1(k0[106]),
        .I2(k0[74]),
        .I3(k0[10]),
        .O(\a1/v3 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair154" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[10]_i_1__0 
       (.I0(k1[42]),
        .I1(k1[106]),
        .I2(k1[74]),
        .I3(k1[10]),
        .O(\a2/v3 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair125" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[10]_i_1__1 
       (.I0(k2[42]),
        .I1(k2[106]),
        .I2(k2[74]),
        .I3(k2[10]),
        .O(\a3/v3 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair92" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[10]_i_1__2 
       (.I0(k3[42]),
        .I1(k3[106]),
        .I2(k3[74]),
        .I3(k3[10]),
        .O(\a4/v3 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair33" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[10]_i_1__3 
       (.I0(k4[42]),
        .I1(k4[106]),
        .I2(k4[74]),
        .I3(k4[10]),
        .O(\a5/v3 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair46" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[10]_i_1__4 
       (.I0(k5[42]),
        .I1(k5[106]),
        .I2(k5[74]),
        .I3(k5[10]),
        .O(\a6/v3 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair271" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[10]_i_1__5 
       (.I0(k6[42]),
        .I1(k6[106]),
        .I2(k6[74]),
        .I3(k6[10]),
        .O(\a7/v3 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair306" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[10]_i_1__6 
       (.I0(k7[42]),
        .I1(k7[106]),
        .I2(k7[74]),
        .I3(k7[10]),
        .O(\a8/v3 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair201" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[10]_i_1__7 
       (.I0(k8[42]),
        .I1(k8[106]),
        .I2(k8[74]),
        .I3(k8[10]),
        .O(\a9/v3 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair233" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[10]_i_1__8 
       (.I0(k9[42]),
        .I1(k9[106]),
        .I2(k9[74]),
        .I3(k9[10]),
        .O(\a10/v3 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair182" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[11]_i_1 
       (.I0(k0[43]),
        .I1(k0[107]),
        .I2(k0[75]),
        .I3(k0[11]),
        .O(\a1/v3 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair153" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[11]_i_1__0 
       (.I0(k1[43]),
        .I1(k1[107]),
        .I2(k1[75]),
        .I3(k1[11]),
        .O(\a2/v3 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair124" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[11]_i_1__1 
       (.I0(k2[43]),
        .I1(k2[107]),
        .I2(k2[75]),
        .I3(k2[11]),
        .O(\a3/v3 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair91" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[11]_i_1__2 
       (.I0(k3[43]),
        .I1(k3[107]),
        .I2(k3[75]),
        .I3(k3[11]),
        .O(\a4/v3 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair32" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[11]_i_1__3 
       (.I0(k4[43]),
        .I1(k4[107]),
        .I2(k4[75]),
        .I3(k4[11]),
        .O(\a5/v3 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair47" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[11]_i_1__4 
       (.I0(k5[43]),
        .I1(k5[107]),
        .I2(k5[75]),
        .I3(k5[11]),
        .O(\a6/v3 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair272" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[11]_i_1__5 
       (.I0(k6[43]),
        .I1(k6[107]),
        .I2(k6[75]),
        .I3(k6[11]),
        .O(\a7/v3 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair305" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[11]_i_1__6 
       (.I0(k7[43]),
        .I1(k7[107]),
        .I2(k7[75]),
        .I3(k7[11]),
        .O(\a8/v3 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair202" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[11]_i_1__7 
       (.I0(k8[43]),
        .I1(k8[107]),
        .I2(k8[75]),
        .I3(k8[11]),
        .O(\a9/v3 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair234" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[11]_i_1__8 
       (.I0(k9[43]),
        .I1(k9[107]),
        .I2(k9[75]),
        .I3(k9[11]),
        .O(\a10/v3 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair181" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[12]_i_1 
       (.I0(k0[44]),
        .I1(k0[108]),
        .I2(k0[76]),
        .I3(k0[12]),
        .O(\a1/v3 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair152" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[12]_i_1__0 
       (.I0(k1[44]),
        .I1(k1[108]),
        .I2(k1[76]),
        .I3(k1[12]),
        .O(\a2/v3 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair123" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[12]_i_1__1 
       (.I0(k2[44]),
        .I1(k2[108]),
        .I2(k2[76]),
        .I3(k2[12]),
        .O(\a3/v3 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[12]_i_1__2 
       (.I0(k3[44]),
        .I1(k3[108]),
        .I2(k3[76]),
        .I3(k3[12]),
        .O(\a4/v3 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair31" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[12]_i_1__3 
       (.I0(k4[44]),
        .I1(k4[108]),
        .I2(k4[76]),
        .I3(k4[12]),
        .O(\a5/v3 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair48" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[12]_i_1__4 
       (.I0(k5[44]),
        .I1(k5[108]),
        .I2(k5[76]),
        .I3(k5[12]),
        .O(\a6/v3 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair273" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[12]_i_1__5 
       (.I0(k6[44]),
        .I1(k6[108]),
        .I2(k6[76]),
        .I3(k6[12]),
        .O(\a7/v3 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair304" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[12]_i_1__6 
       (.I0(k7[44]),
        .I1(k7[108]),
        .I2(k7[76]),
        .I3(k7[12]),
        .O(\a8/v3 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair203" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[12]_i_1__7 
       (.I0(k8[44]),
        .I1(k8[108]),
        .I2(k8[76]),
        .I3(k8[12]),
        .O(\a9/v3 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair235" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[12]_i_1__8 
       (.I0(k9[44]),
        .I1(k9[108]),
        .I2(k9[76]),
        .I3(k9[12]),
        .O(\a10/v3 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair180" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[13]_i_1 
       (.I0(k0[45]),
        .I1(k0[109]),
        .I2(k0[77]),
        .I3(k0[13]),
        .O(\a1/v3 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair151" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[13]_i_1__0 
       (.I0(k1[45]),
        .I1(k1[109]),
        .I2(k1[77]),
        .I3(k1[13]),
        .O(\a2/v3 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair122" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[13]_i_1__1 
       (.I0(k2[45]),
        .I1(k2[109]),
        .I2(k2[77]),
        .I3(k2[13]),
        .O(\a3/v3 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair89" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[13]_i_1__2 
       (.I0(k3[45]),
        .I1(k3[109]),
        .I2(k3[77]),
        .I3(k3[13]),
        .O(\a4/v3 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair30" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[13]_i_1__3 
       (.I0(k4[45]),
        .I1(k4[109]),
        .I2(k4[77]),
        .I3(k4[13]),
        .O(\a5/v3 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair49" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[13]_i_1__4 
       (.I0(k5[45]),
        .I1(k5[109]),
        .I2(k5[77]),
        .I3(k5[13]),
        .O(\a6/v3 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair274" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[13]_i_1__5 
       (.I0(k6[45]),
        .I1(k6[109]),
        .I2(k6[77]),
        .I3(k6[13]),
        .O(\a7/v3 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair303" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[13]_i_1__6 
       (.I0(k7[45]),
        .I1(k7[109]),
        .I2(k7[77]),
        .I3(k7[13]),
        .O(\a8/v3 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair204" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[13]_i_1__7 
       (.I0(k8[45]),
        .I1(k8[109]),
        .I2(k8[77]),
        .I3(k8[13]),
        .O(\a9/v3 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair236" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[13]_i_1__8 
       (.I0(k9[45]),
        .I1(k9[109]),
        .I2(k9[77]),
        .I3(k9[13]),
        .O(\a10/v3 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair179" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[14]_i_1 
       (.I0(k0[46]),
        .I1(k0[110]),
        .I2(k0[78]),
        .I3(k0[14]),
        .O(\a1/v3 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair150" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[14]_i_1__0 
       (.I0(k1[46]),
        .I1(k1[110]),
        .I2(k1[78]),
        .I3(k1[14]),
        .O(\a2/v3 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair121" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[14]_i_1__1 
       (.I0(k2[46]),
        .I1(k2[110]),
        .I2(k2[78]),
        .I3(k2[14]),
        .O(\a3/v3 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair88" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[14]_i_1__2 
       (.I0(k3[46]),
        .I1(k3[110]),
        .I2(k3[78]),
        .I3(k3[14]),
        .O(\a4/v3 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair29" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[14]_i_1__3 
       (.I0(k4[46]),
        .I1(k4[110]),
        .I2(k4[78]),
        .I3(k4[14]),
        .O(\a5/v3 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair50" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[14]_i_1__4 
       (.I0(k5[46]),
        .I1(k5[110]),
        .I2(k5[78]),
        .I3(k5[14]),
        .O(\a6/v3 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair275" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[14]_i_1__5 
       (.I0(k6[46]),
        .I1(k6[110]),
        .I2(k6[78]),
        .I3(k6[14]),
        .O(\a7/v3 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair302" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[14]_i_1__6 
       (.I0(k7[46]),
        .I1(k7[110]),
        .I2(k7[78]),
        .I3(k7[14]),
        .O(\a8/v3 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair205" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[14]_i_1__7 
       (.I0(k8[46]),
        .I1(k8[110]),
        .I2(k8[78]),
        .I3(k8[14]),
        .O(\a9/v3 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair237" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[14]_i_1__8 
       (.I0(k9[46]),
        .I1(k9[110]),
        .I2(k9[78]),
        .I3(k9[14]),
        .O(\a10/v3 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair178" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[15]_i_1 
       (.I0(k0[47]),
        .I1(k0[111]),
        .I2(k0[79]),
        .I3(k0[15]),
        .O(\a1/v3 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair149" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[15]_i_1__0 
       (.I0(k1[47]),
        .I1(k1[111]),
        .I2(k1[79]),
        .I3(k1[15]),
        .O(\a2/v3 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair120" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[15]_i_1__1 
       (.I0(k2[47]),
        .I1(k2[111]),
        .I2(k2[79]),
        .I3(k2[15]),
        .O(\a3/v3 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair87" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[15]_i_1__2 
       (.I0(k3[47]),
        .I1(k3[111]),
        .I2(k3[79]),
        .I3(k3[15]),
        .O(\a4/v3 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair28" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[15]_i_1__3 
       (.I0(k4[47]),
        .I1(k4[111]),
        .I2(k4[79]),
        .I3(k4[15]),
        .O(\a5/v3 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair51" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[15]_i_1__4 
       (.I0(k5[47]),
        .I1(k5[111]),
        .I2(k5[79]),
        .I3(k5[15]),
        .O(\a6/v3 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair276" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[15]_i_1__5 
       (.I0(k6[47]),
        .I1(k6[111]),
        .I2(k6[79]),
        .I3(k6[15]),
        .O(\a7/v3 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair301" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[15]_i_1__6 
       (.I0(k7[47]),
        .I1(k7[111]),
        .I2(k7[79]),
        .I3(k7[15]),
        .O(\a8/v3 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair206" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[15]_i_1__7 
       (.I0(k8[47]),
        .I1(k8[111]),
        .I2(k8[79]),
        .I3(k8[15]),
        .O(\a9/v3 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair238" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[15]_i_1__8 
       (.I0(k9[47]),
        .I1(k9[111]),
        .I2(k9[79]),
        .I3(k9[15]),
        .O(\a10/v3 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair177" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[16]_i_1 
       (.I0(k0[48]),
        .I1(k0[112]),
        .I2(k0[80]),
        .I3(k0[16]),
        .O(\a1/v3 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair148" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[16]_i_1__0 
       (.I0(k1[48]),
        .I1(k1[112]),
        .I2(k1[80]),
        .I3(k1[16]),
        .O(\a2/v3 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair119" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[16]_i_1__1 
       (.I0(k2[48]),
        .I1(k2[112]),
        .I2(k2[80]),
        .I3(k2[16]),
        .O(\a3/v3 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair86" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[16]_i_1__2 
       (.I0(k3[48]),
        .I1(k3[112]),
        .I2(k3[80]),
        .I3(k3[16]),
        .O(\a4/v3 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair27" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[16]_i_1__3 
       (.I0(k4[48]),
        .I1(k4[112]),
        .I2(k4[80]),
        .I3(k4[16]),
        .O(\a5/v3 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair52" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[16]_i_1__4 
       (.I0(k5[48]),
        .I1(k5[112]),
        .I2(k5[80]),
        .I3(k5[16]),
        .O(\a6/v3 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair277" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[16]_i_1__5 
       (.I0(k6[48]),
        .I1(k6[112]),
        .I2(k6[80]),
        .I3(k6[16]),
        .O(\a7/v3 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair300" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[16]_i_1__6 
       (.I0(k7[48]),
        .I1(k7[112]),
        .I2(k7[80]),
        .I3(k7[16]),
        .O(\a8/v3 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair207" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[16]_i_1__7 
       (.I0(k8[48]),
        .I1(k8[112]),
        .I2(k8[80]),
        .I3(k8[16]),
        .O(\a9/v3 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair239" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[16]_i_1__8 
       (.I0(k9[48]),
        .I1(k9[112]),
        .I2(k9[80]),
        .I3(k9[16]),
        .O(\a10/v3 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair176" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[17]_i_1 
       (.I0(k0[49]),
        .I1(k0[113]),
        .I2(k0[81]),
        .I3(k0[17]),
        .O(\a1/v3 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair147" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[17]_i_1__0 
       (.I0(k1[49]),
        .I1(k1[113]),
        .I2(k1[81]),
        .I3(k1[17]),
        .O(\a2/v3 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair118" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[17]_i_1__1 
       (.I0(k2[49]),
        .I1(k2[113]),
        .I2(k2[81]),
        .I3(k2[17]),
        .O(\a3/v3 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair85" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[17]_i_1__2 
       (.I0(k3[49]),
        .I1(k3[113]),
        .I2(k3[81]),
        .I3(k3[17]),
        .O(\a4/v3 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair102" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[17]_i_1__3 
       (.I0(k4[49]),
        .I1(k4[113]),
        .I2(k4[81]),
        .I3(k4[17]),
        .O(\a5/v3 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair53" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[17]_i_1__4 
       (.I0(k5[49]),
        .I1(k5[113]),
        .I2(k5[81]),
        .I3(k5[17]),
        .O(\a6/v3 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair278" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[17]_i_1__5 
       (.I0(k6[49]),
        .I1(k6[113]),
        .I2(k6[81]),
        .I3(k6[17]),
        .O(\a7/v3 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair299" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[17]_i_1__6 
       (.I0(k7[49]),
        .I1(k7[113]),
        .I2(k7[81]),
        .I3(k7[17]),
        .O(\a8/v3 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair208" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[17]_i_1__7 
       (.I0(k8[49]),
        .I1(k8[113]),
        .I2(k8[81]),
        .I3(k8[17]),
        .O(\a9/v3 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair240" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[17]_i_1__8 
       (.I0(k9[49]),
        .I1(k9[113]),
        .I2(k9[81]),
        .I3(k9[17]),
        .O(\a10/v3 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair175" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[18]_i_1 
       (.I0(k0[50]),
        .I1(k0[114]),
        .I2(k0[82]),
        .I3(k0[18]),
        .O(\a1/v3 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair146" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[18]_i_1__0 
       (.I0(k1[50]),
        .I1(k1[114]),
        .I2(k1[82]),
        .I3(k1[18]),
        .O(\a2/v3 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair117" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[18]_i_1__1 
       (.I0(k2[50]),
        .I1(k2[114]),
        .I2(k2[82]),
        .I3(k2[18]),
        .O(\a3/v3 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair84" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[18]_i_1__2 
       (.I0(k3[50]),
        .I1(k3[114]),
        .I2(k3[82]),
        .I3(k3[18]),
        .O(\a4/v3 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair25" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[18]_i_1__3 
       (.I0(k4[50]),
        .I1(k4[114]),
        .I2(k4[82]),
        .I3(k4[18]),
        .O(\a5/v3 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair54" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[18]_i_1__4 
       (.I0(k5[50]),
        .I1(k5[114]),
        .I2(k5[82]),
        .I3(k5[18]),
        .O(\a6/v3 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair279" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[18]_i_1__5 
       (.I0(k6[50]),
        .I1(k6[114]),
        .I2(k6[82]),
        .I3(k6[18]),
        .O(\a7/v3 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair298" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[18]_i_1__6 
       (.I0(k7[50]),
        .I1(k7[114]),
        .I2(k7[82]),
        .I3(k7[18]),
        .O(\a8/v3 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair209" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[18]_i_1__7 
       (.I0(k8[50]),
        .I1(k8[114]),
        .I2(k8[82]),
        .I3(k8[18]),
        .O(\a9/v3 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair241" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[18]_i_1__8 
       (.I0(k9[50]),
        .I1(k9[114]),
        .I2(k9[82]),
        .I3(k9[18]),
        .O(\a10/v3 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair174" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[19]_i_1 
       (.I0(k0[51]),
        .I1(k0[115]),
        .I2(k0[83]),
        .I3(k0[19]),
        .O(\a1/v3 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair145" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[19]_i_1__0 
       (.I0(k1[51]),
        .I1(k1[115]),
        .I2(k1[83]),
        .I3(k1[19]),
        .O(\a2/v3 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair116" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[19]_i_1__1 
       (.I0(k2[51]),
        .I1(k2[115]),
        .I2(k2[83]),
        .I3(k2[19]),
        .O(\a3/v3 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair83" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[19]_i_1__2 
       (.I0(k3[51]),
        .I1(k3[115]),
        .I2(k3[83]),
        .I3(k3[19]),
        .O(\a4/v3 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair24" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[19]_i_1__3 
       (.I0(k4[51]),
        .I1(k4[115]),
        .I2(k4[83]),
        .I3(k4[19]),
        .O(\a5/v3 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair55" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[19]_i_1__4 
       (.I0(k5[51]),
        .I1(k5[115]),
        .I2(k5[83]),
        .I3(k5[19]),
        .O(\a6/v3 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair280" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[19]_i_1__5 
       (.I0(k6[51]),
        .I1(k6[115]),
        .I2(k6[83]),
        .I3(k6[19]),
        .O(\a7/v3 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair297" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[19]_i_1__6 
       (.I0(k7[51]),
        .I1(k7[115]),
        .I2(k7[83]),
        .I3(k7[19]),
        .O(\a8/v3 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair210" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[19]_i_1__7 
       (.I0(k8[51]),
        .I1(k8[115]),
        .I2(k8[83]),
        .I3(k8[19]),
        .O(\a9/v3 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair242" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[19]_i_1__8 
       (.I0(k9[51]),
        .I1(k9[115]),
        .I2(k9[83]),
        .I3(k9[19]),
        .O(\a10/v3 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair103" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[1]_i_1 
       (.I0(k0[33]),
        .I1(k0[97]),
        .I2(k0[65]),
        .I3(k0[1]),
        .O(\a1/v3 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair11" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[1]_i_1__0 
       (.I0(k1[33]),
        .I1(k1[97]),
        .I2(k1[65]),
        .I3(k1[1]),
        .O(\a2/v3 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair10" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[1]_i_1__1 
       (.I0(k2[33]),
        .I1(k2[97]),
        .I2(k2[65]),
        .I3(k2[1]),
        .O(\a3/v3 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[1]_i_1__2 
       (.I0(k3[33]),
        .I1(k3[97]),
        .I2(k3[65]),
        .I3(k3[1]),
        .O(\a4/v3 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[1]_i_1__3 
       (.I0(k4[33]),
        .I1(k4[97]),
        .I2(k4[65]),
        .I3(k4[1]),
        .O(\a5/v3 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair37" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[1]_i_1__4 
       (.I0(k5[33]),
        .I1(k5[97]),
        .I2(k5[65]),
        .I3(k5[1]),
        .O(\a6/v3 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair262" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[1]_i_1__5 
       (.I0(k6[33]),
        .I1(k6[97]),
        .I2(k6[65]),
        .I3(k6[1]),
        .O(\a7/v3 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair315" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[1]_i_1__6 
       (.I0(k7[33]),
        .I1(k7[97]),
        .I2(k7[65]),
        .I3(k7[1]),
        .O(\a8/v3 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair318" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[1]_i_1__7 
       (.I0(k8[33]),
        .I1(k8[97]),
        .I2(k8[65]),
        .I3(k8[1]),
        .O(\a9/v3 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair224" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[1]_i_1__8 
       (.I0(k9[33]),
        .I1(k9[97]),
        .I2(k9[65]),
        .I3(k9[1]),
        .O(\a10/v3 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair173" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[20]_i_1 
       (.I0(k0[52]),
        .I1(k0[116]),
        .I2(k0[84]),
        .I3(k0[20]),
        .O(\a1/v3 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair144" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[20]_i_1__0 
       (.I0(k1[52]),
        .I1(k1[116]),
        .I2(k1[84]),
        .I3(k1[20]),
        .O(\a2/v3 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair115" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[20]_i_1__1 
       (.I0(k2[52]),
        .I1(k2[116]),
        .I2(k2[84]),
        .I3(k2[20]),
        .O(\a3/v3 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair82" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[20]_i_1__2 
       (.I0(k3[52]),
        .I1(k3[116]),
        .I2(k3[84]),
        .I3(k3[20]),
        .O(\a4/v3 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair23" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[20]_i_1__3 
       (.I0(k4[52]),
        .I1(k4[116]),
        .I2(k4[84]),
        .I3(k4[20]),
        .O(\a5/v3 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair56" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[20]_i_1__4 
       (.I0(k5[52]),
        .I1(k5[116]),
        .I2(k5[84]),
        .I3(k5[20]),
        .O(\a6/v3 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair281" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[20]_i_1__5 
       (.I0(k6[52]),
        .I1(k6[116]),
        .I2(k6[84]),
        .I3(k6[20]),
        .O(\a7/v3 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair296" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[20]_i_1__6 
       (.I0(k7[52]),
        .I1(k7[116]),
        .I2(k7[84]),
        .I3(k7[20]),
        .O(\a8/v3 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair211" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[20]_i_1__7 
       (.I0(k8[52]),
        .I1(k8[116]),
        .I2(k8[84]),
        .I3(k8[20]),
        .O(\a9/v3 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair243" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[20]_i_1__8 
       (.I0(k9[52]),
        .I1(k9[116]),
        .I2(k9[84]),
        .I3(k9[20]),
        .O(\a10/v3 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair172" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[21]_i_1 
       (.I0(k0[53]),
        .I1(k0[117]),
        .I2(k0[85]),
        .I3(k0[21]),
        .O(\a1/v3 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair143" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[21]_i_1__0 
       (.I0(k1[53]),
        .I1(k1[117]),
        .I2(k1[85]),
        .I3(k1[21]),
        .O(\a2/v3 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair114" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[21]_i_1__1 
       (.I0(k2[53]),
        .I1(k2[117]),
        .I2(k2[85]),
        .I3(k2[21]),
        .O(\a3/v3 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair81" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[21]_i_1__2 
       (.I0(k3[53]),
        .I1(k3[117]),
        .I2(k3[85]),
        .I3(k3[21]),
        .O(\a4/v3 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair22" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[21]_i_1__3 
       (.I0(k4[53]),
        .I1(k4[117]),
        .I2(k4[85]),
        .I3(k4[21]),
        .O(\a5/v3 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair57" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[21]_i_1__4 
       (.I0(k5[53]),
        .I1(k5[117]),
        .I2(k5[85]),
        .I3(k5[21]),
        .O(\a6/v3 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair282" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[21]_i_1__5 
       (.I0(k6[53]),
        .I1(k6[117]),
        .I2(k6[85]),
        .I3(k6[21]),
        .O(\a7/v3 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair295" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[21]_i_1__6 
       (.I0(k7[53]),
        .I1(k7[117]),
        .I2(k7[85]),
        .I3(k7[21]),
        .O(\a8/v3 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair212" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[21]_i_1__7 
       (.I0(k8[53]),
        .I1(k8[117]),
        .I2(k8[85]),
        .I3(k8[21]),
        .O(\a9/v3 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair244" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[21]_i_1__8 
       (.I0(k9[53]),
        .I1(k9[117]),
        .I2(k9[85]),
        .I3(k9[21]),
        .O(\a10/v3 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair171" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[22]_i_1 
       (.I0(k0[54]),
        .I1(k0[118]),
        .I2(k0[86]),
        .I3(k0[22]),
        .O(\a1/v3 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair142" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[22]_i_1__0 
       (.I0(k1[54]),
        .I1(k1[118]),
        .I2(k1[86]),
        .I3(k1[22]),
        .O(\a2/v3 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair113" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[22]_i_1__1 
       (.I0(k2[54]),
        .I1(k2[118]),
        .I2(k2[86]),
        .I3(k2[22]),
        .O(\a3/v3 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair80" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[22]_i_1__2 
       (.I0(k3[54]),
        .I1(k3[118]),
        .I2(k3[86]),
        .I3(k3[22]),
        .O(\a4/v3 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair21" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[22]_i_1__3 
       (.I0(k4[54]),
        .I1(k4[118]),
        .I2(k4[86]),
        .I3(k4[22]),
        .O(\a5/v3 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair58" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[22]_i_1__4 
       (.I0(k5[54]),
        .I1(k5[118]),
        .I2(k5[86]),
        .I3(k5[22]),
        .O(\a6/v3 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair283" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[22]_i_1__5 
       (.I0(k6[54]),
        .I1(k6[118]),
        .I2(k6[86]),
        .I3(k6[22]),
        .O(\a7/v3 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair294" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[22]_i_1__6 
       (.I0(k7[54]),
        .I1(k7[118]),
        .I2(k7[86]),
        .I3(k7[22]),
        .O(\a8/v3 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair213" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[22]_i_1__7 
       (.I0(k8[54]),
        .I1(k8[118]),
        .I2(k8[86]),
        .I3(k8[22]),
        .O(\a9/v3 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair245" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[22]_i_1__8 
       (.I0(k9[54]),
        .I1(k9[118]),
        .I2(k9[86]),
        .I3(k9[22]),
        .O(\a10/v3 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair170" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[23]_i_1 
       (.I0(k0[55]),
        .I1(k0[119]),
        .I2(k0[87]),
        .I3(k0[23]),
        .O(\a1/v3 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair141" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[23]_i_1__0 
       (.I0(k1[55]),
        .I1(k1[119]),
        .I2(k1[87]),
        .I3(k1[23]),
        .O(\a2/v3 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair112" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[23]_i_1__1 
       (.I0(k2[55]),
        .I1(k2[119]),
        .I2(k2[87]),
        .I3(k2[23]),
        .O(\a3/v3 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair79" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[23]_i_1__2 
       (.I0(k3[55]),
        .I1(k3[119]),
        .I2(k3[87]),
        .I3(k3[23]),
        .O(\a4/v3 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair20" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[23]_i_1__3 
       (.I0(k4[55]),
        .I1(k4[119]),
        .I2(k4[87]),
        .I3(k4[23]),
        .O(\a5/v3 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair59" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[23]_i_1__4 
       (.I0(k5[55]),
        .I1(k5[119]),
        .I2(k5[87]),
        .I3(k5[23]),
        .O(\a6/v3 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair284" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[23]_i_1__5 
       (.I0(k6[55]),
        .I1(k6[119]),
        .I2(k6[87]),
        .I3(k6[23]),
        .O(\a7/v3 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair317" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[23]_i_1__6 
       (.I0(k7[55]),
        .I1(k7[119]),
        .I2(k7[87]),
        .I3(k7[23]),
        .O(\a8/v3 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair214" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[23]_i_1__7 
       (.I0(k8[55]),
        .I1(k8[119]),
        .I2(k8[87]),
        .I3(k8[23]),
        .O(\a9/v3 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair246" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[23]_i_1__8 
       (.I0(k9[55]),
        .I1(k9[119]),
        .I2(k9[87]),
        .I3(k9[23]),
        .O(\a10/v3 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair162" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    \k3a[24]_i_1 
       (.I0(k0[56]),
        .I1(k0[120]),
        .I2(k0[88]),
        .I3(k0[24]),
        .O(\a1/v3 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair140" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[24]_i_1__0 
       (.I0(k1[56]),
        .I1(k1[120]),
        .I2(k1[88]),
        .I3(k1[24]),
        .O(\a2/v3 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair111" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[24]_i_1__1 
       (.I0(k2[56]),
        .I1(k2[120]),
        .I2(k2[88]),
        .I3(k2[24]),
        .O(\a3/v3 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair78" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[24]_i_1__2 
       (.I0(k3[56]),
        .I1(k3[120]),
        .I2(k3[88]),
        .I3(k3[24]),
        .O(\a4/v3 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair19" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[24]_i_1__3 
       (.I0(k4[56]),
        .I1(k4[120]),
        .I2(k4[88]),
        .I3(k4[24]),
        .O(\a5/v3 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair60" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[24]_i_1__4 
       (.I0(k5[56]),
        .I1(k5[120]),
        .I2(k5[88]),
        .I3(k5[24]),
        .O(\a6/v3 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair285" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[24]_i_1__5 
       (.I0(k6[56]),
        .I1(k6[120]),
        .I2(k6[88]),
        .I3(k6[24]),
        .O(\a7/v3 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair260" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[24]_i_1__6 
       (.I0(k7[56]),
        .I1(k7[120]),
        .I2(k7[88]),
        .I3(k7[24]),
        .O(\a8/v3 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair219" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    \k3a[24]_i_1__7 
       (.I0(k8[56]),
        .I1(k8[120]),
        .I2(k8[88]),
        .I3(k8[24]),
        .O(\a9/v3 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair247" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[24]_i_1__8 
       (.I0(k9[56]),
        .I1(k9[120]),
        .I2(k9[88]),
        .I3(k9[24]),
        .O(\a10/v3 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair169" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[25]_i_1 
       (.I0(k0[57]),
        .I1(k0[121]),
        .I2(k0[89]),
        .I3(k0[25]),
        .O(\a1/v3 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair133" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    \k3a[25]_i_1__0 
       (.I0(k1[57]),
        .I1(k1[121]),
        .I2(k1[89]),
        .I3(k1[25]),
        .O(\a2/v3 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair110" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[25]_i_1__1 
       (.I0(k2[57]),
        .I1(k2[121]),
        .I2(k2[89]),
        .I3(k2[25]),
        .O(\a3/v3 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair77" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[25]_i_1__2 
       (.I0(k3[57]),
        .I1(k3[121]),
        .I2(k3[89]),
        .I3(k3[25]),
        .O(\a4/v3 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair18" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[25]_i_1__3 
       (.I0(k4[57]),
        .I1(k4[121]),
        .I2(k4[89]),
        .I3(k4[25]),
        .O(\a5/v3 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair61" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[25]_i_1__4 
       (.I0(k5[57]),
        .I1(k5[121]),
        .I2(k5[89]),
        .I3(k5[25]),
        .O(\a6/v3 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair286" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[25]_i_1__5 
       (.I0(k6[57]),
        .I1(k6[121]),
        .I2(k6[89]),
        .I3(k6[25]),
        .O(\a7/v3 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair259" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[25]_i_1__6 
       (.I0(k7[57]),
        .I1(k7[121]),
        .I2(k7[89]),
        .I3(k7[25]),
        .O(\a8/v3 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair220" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    \k3a[25]_i_1__7 
       (.I0(k8[57]),
        .I1(k8[121]),
        .I2(k8[89]),
        .I3(k8[25]),
        .O(\a9/v3 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair251" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    \k3a[25]_i_1__8 
       (.I0(k9[57]),
        .I1(k9[121]),
        .I2(k9[89]),
        .I3(k9[25]),
        .O(\a10/v3 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair168" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[26]_i_1 
       (.I0(k0[58]),
        .I1(k0[122]),
        .I2(k0[90]),
        .I3(k0[26]),
        .O(\a1/v3 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair139" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[26]_i_1__0 
       (.I0(k1[58]),
        .I1(k1[122]),
        .I2(k1[90]),
        .I3(k1[26]),
        .O(\a2/v3 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair104" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    \k3a[26]_i_1__1 
       (.I0(k2[58]),
        .I1(k2[122]),
        .I2(k2[90]),
        .I3(k2[26]),
        .O(\a3/v3 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair76" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[26]_i_1__2 
       (.I0(k3[58]),
        .I1(k3[122]),
        .I2(k3[90]),
        .I3(k3[26]),
        .O(\a4/v3 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair17" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[26]_i_1__3 
       (.I0(k4[58]),
        .I1(k4[122]),
        .I2(k4[90]),
        .I3(k4[26]),
        .O(\a5/v3 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair62" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[26]_i_1__4 
       (.I0(k5[58]),
        .I1(k5[122]),
        .I2(k5[90]),
        .I3(k5[26]),
        .O(\a6/v3 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair287" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[26]_i_1__5 
       (.I0(k6[58]),
        .I1(k6[122]),
        .I2(k6[90]),
        .I3(k6[26]),
        .O(\a7/v3 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair258" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[26]_i_1__6 
       (.I0(k7[58]),
        .I1(k7[122]),
        .I2(k7[90]),
        .I3(k7[26]),
        .O(\a8/v3 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair215" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[26]_i_1__7 
       (.I0(k8[58]),
        .I1(k8[122]),
        .I2(k8[90]),
        .I3(k8[26]),
        .O(\a9/v3 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair252" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    \k3a[26]_i_1__8 
       (.I0(k9[58]),
        .I1(k9[122]),
        .I2(k9[90]),
        .I3(k9[26]),
        .O(\a10/v3 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair167" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[27]_i_1 
       (.I0(k0[59]),
        .I1(k0[123]),
        .I2(k0[91]),
        .I3(k0[27]),
        .O(\a1/v3 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair138" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[27]_i_1__0 
       (.I0(k1[59]),
        .I1(k1[123]),
        .I2(k1[91]),
        .I3(k1[27]),
        .O(\a2/v3 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair109" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[27]_i_1__1 
       (.I0(k2[59]),
        .I1(k2[123]),
        .I2(k2[91]),
        .I3(k2[27]),
        .O(\a3/v3 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair71" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    \k3a[27]_i_1__2 
       (.I0(k3[59]),
        .I1(k3[123]),
        .I2(k3[91]),
        .I3(k3[27]),
        .O(\a4/v3 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair16" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[27]_i_1__3 
       (.I0(k4[59]),
        .I1(k4[123]),
        .I2(k4[91]),
        .I3(k4[27]),
        .O(\a5/v3 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair63" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[27]_i_1__4 
       (.I0(k5[59]),
        .I1(k5[123]),
        .I2(k5[91]),
        .I3(k5[27]),
        .O(\a6/v3 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair288" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[27]_i_1__5 
       (.I0(k6[59]),
        .I1(k6[123]),
        .I2(k6[91]),
        .I3(k6[27]),
        .O(\a7/v3 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair257" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[27]_i_1__6 
       (.I0(k7[59]),
        .I1(k7[123]),
        .I2(k7[91]),
        .I3(k7[27]),
        .O(\a8/v3 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair221" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    \k3a[27]_i_1__7 
       (.I0(k8[59]),
        .I1(k8[123]),
        .I2(k8[91]),
        .I3(k8[27]),
        .O(\a9/v3 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair248" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[27]_i_1__8 
       (.I0(k9[59]),
        .I1(k9[123]),
        .I2(k9[91]),
        .I3(k9[27]),
        .O(\a10/v3 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair166" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[28]_i_1 
       (.I0(k0[60]),
        .I1(k0[124]),
        .I2(k0[92]),
        .I3(k0[28]),
        .O(\a1/v3 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair137" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[28]_i_1__0 
       (.I0(k1[60]),
        .I1(k1[124]),
        .I2(k1[92]),
        .I3(k1[28]),
        .O(\a2/v3 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair108" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[28]_i_1__1 
       (.I0(k2[60]),
        .I1(k2[124]),
        .I2(k2[92]),
        .I3(k2[28]),
        .O(\a3/v3 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair75" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[28]_i_1__2 
       (.I0(k3[60]),
        .I1(k3[124]),
        .I2(k3[92]),
        .I3(k3[28]),
        .O(\a4/v3 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair12" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    \k3a[28]_i_1__3 
       (.I0(k4[60]),
        .I1(k4[124]),
        .I2(k4[92]),
        .I3(k4[28]),
        .O(\a5/v3 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair64" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[28]_i_1__4 
       (.I0(k5[60]),
        .I1(k5[124]),
        .I2(k5[92]),
        .I3(k5[28]),
        .O(\a6/v3 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair289" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[28]_i_1__5 
       (.I0(k6[60]),
        .I1(k6[124]),
        .I2(k6[92]),
        .I3(k6[28]),
        .O(\a7/v3 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair256" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[28]_i_1__6 
       (.I0(k7[60]),
        .I1(k7[124]),
        .I2(k7[92]),
        .I3(k7[28]),
        .O(\a8/v3 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair222" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    \k3a[28]_i_1__7 
       (.I0(k8[60]),
        .I1(k8[124]),
        .I2(k8[92]),
        .I3(k8[28]),
        .O(\a9/v3 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair253" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    \k3a[28]_i_1__8 
       (.I0(k9[60]),
        .I1(k9[124]),
        .I2(k9[92]),
        .I3(k9[28]),
        .O(\a10/v3 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair165" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[29]_i_1 
       (.I0(k0[61]),
        .I1(k0[125]),
        .I2(k0[93]),
        .I3(k0[29]),
        .O(\a1/v3 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair136" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[29]_i_1__0 
       (.I0(k1[61]),
        .I1(k1[125]),
        .I2(k1[93]),
        .I3(k1[29]),
        .O(\a2/v3 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair107" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[29]_i_1__1 
       (.I0(k2[61]),
        .I1(k2[125]),
        .I2(k2[93]),
        .I3(k2[29]),
        .O(\a3/v3 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair74" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[29]_i_1__2 
       (.I0(k3[61]),
        .I1(k3[125]),
        .I2(k3[93]),
        .I3(k3[29]),
        .O(\a4/v3 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair15" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[29]_i_1__3 
       (.I0(k4[61]),
        .I1(k4[125]),
        .I2(k4[93]),
        .I3(k4[29]),
        .O(\a5/v3 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair67" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    \k3a[29]_i_1__4 
       (.I0(k5[61]),
        .I1(k5[125]),
        .I2(k5[93]),
        .I3(k5[29]),
        .O(\a6/v3 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair290" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[29]_i_1__5 
       (.I0(k6[61]),
        .I1(k6[125]),
        .I2(k6[93]),
        .I3(k6[29]),
        .O(\a7/v3 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair255" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[29]_i_1__6 
       (.I0(k7[61]),
        .I1(k7[125]),
        .I2(k7[93]),
        .I3(k7[29]),
        .O(\a8/v3 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair216" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[29]_i_1__7 
       (.I0(k8[61]),
        .I1(k8[125]),
        .I2(k8[93]),
        .I3(k8[29]),
        .O(\a9/v3 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair254" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    \k3a[29]_i_1__8 
       (.I0(k9[61]),
        .I1(k9[125]),
        .I2(k9[93]),
        .I3(k9[29]),
        .O(\a10/v3 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair191" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[2]_i_1 
       (.I0(k0[34]),
        .I1(k0[98]),
        .I2(k0[66]),
        .I3(k0[2]),
        .O(\a1/v3 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[2]_i_1__0 
       (.I0(k1[34]),
        .I1(k1[98]),
        .I2(k1[66]),
        .I3(k1[2]),
        .O(\a2/v3 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[2]_i_1__1 
       (.I0(k2[34]),
        .I1(k2[98]),
        .I2(k2[66]),
        .I3(k2[2]),
        .O(\a3/v3 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair100" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[2]_i_1__2 
       (.I0(k3[34]),
        .I1(k3[98]),
        .I2(k3[66]),
        .I3(k3[2]),
        .O(\a4/v3 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair35" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[2]_i_1__3 
       (.I0(k4[34]),
        .I1(k4[98]),
        .I2(k4[66]),
        .I3(k4[2]),
        .O(\a5/v3 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair38" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[2]_i_1__4 
       (.I0(k5[34]),
        .I1(k5[98]),
        .I2(k5[66]),
        .I3(k5[2]),
        .O(\a6/v3 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair263" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[2]_i_1__5 
       (.I0(k6[34]),
        .I1(k6[98]),
        .I2(k6[66]),
        .I3(k6[2]),
        .O(\a7/v3 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair314" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[2]_i_1__6 
       (.I0(k7[34]),
        .I1(k7[98]),
        .I2(k7[66]),
        .I3(k7[2]),
        .O(\a8/v3 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair193" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[2]_i_1__7 
       (.I0(k8[34]),
        .I1(k8[98]),
        .I2(k8[66]),
        .I3(k8[2]),
        .O(\a9/v3 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair225" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[2]_i_1__8 
       (.I0(k9[34]),
        .I1(k9[98]),
        .I2(k9[66]),
        .I3(k9[2]),
        .O(\a10/v3 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair164" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[30]_i_1 
       (.I0(k0[62]),
        .I1(k0[126]),
        .I2(k0[94]),
        .I3(k0[30]),
        .O(\a1/v3 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair135" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[30]_i_1__0 
       (.I0(k1[62]),
        .I1(k1[126]),
        .I2(k1[94]),
        .I3(k1[30]),
        .O(\a2/v3 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair106" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[30]_i_1__1 
       (.I0(k2[62]),
        .I1(k2[126]),
        .I2(k2[94]),
        .I3(k2[30]),
        .O(\a3/v3 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair73" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[30]_i_1__2 
       (.I0(k3[62]),
        .I1(k3[126]),
        .I2(k3[94]),
        .I3(k3[30]),
        .O(\a4/v3 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[30]_i_1__3 
       (.I0(k4[62]),
        .I1(k4[126]),
        .I2(k4[94]),
        .I3(k4[30]),
        .O(\a5/v3 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair65" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[30]_i_1__4 
       (.I0(k5[62]),
        .I1(k5[126]),
        .I2(k5[94]),
        .I3(k5[30]),
        .O(\a6/v3 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair292" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    \k3a[30]_i_1__5 
       (.I0(k6[62]),
        .I1(k6[126]),
        .I2(k6[94]),
        .I3(k6[30]),
        .O(\a7/v3 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair293" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[30]_i_1__6 
       (.I0(k7[62]),
        .I1(k7[126]),
        .I2(k7[94]),
        .I3(k7[30]),
        .O(\a8/v3 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair217" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[30]_i_1__7 
       (.I0(k8[62]),
        .I1(k8[126]),
        .I2(k8[94]),
        .I3(k8[30]),
        .O(\a9/v3 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair249" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[30]_i_1__8 
       (.I0(k9[62]),
        .I1(k9[126]),
        .I2(k9[94]),
        .I3(k9[30]),
        .O(\a10/v3 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair163" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[31]_i_1 
       (.I0(k0[63]),
        .I1(k0[127]),
        .I2(k0[95]),
        .I3(k0[31]),
        .O(\a1/v3 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair134" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[31]_i_1__0 
       (.I0(k1[63]),
        .I1(k1[127]),
        .I2(k1[95]),
        .I3(k1[31]),
        .O(\a2/v3 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair105" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[31]_i_1__1 
       (.I0(k2[63]),
        .I1(k2[127]),
        .I2(k2[95]),
        .I3(k2[31]),
        .O(\a3/v3 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair72" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[31]_i_1__2 
       (.I0(k3[63]),
        .I1(k3[127]),
        .I2(k3[95]),
        .I3(k3[31]),
        .O(\a4/v3 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[31]_i_1__3 
       (.I0(k4[63]),
        .I1(k4[127]),
        .I2(k4[95]),
        .I3(k4[31]),
        .O(\a5/v3 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair66" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[31]_i_1__4 
       (.I0(k5[63]),
        .I1(k5[127]),
        .I2(k5[95]),
        .I3(k5[31]),
        .O(\a6/v3 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair291" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[31]_i_1__5 
       (.I0(k6[63]),
        .I1(k6[127]),
        .I2(k6[95]),
        .I3(k6[31]),
        .O(\a7/v3 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair319" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    \k3a[31]_i_1__6 
       (.I0(k7[63]),
        .I1(k7[127]),
        .I2(k7[95]),
        .I3(k7[31]),
        .O(\a8/v3 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair218" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[31]_i_1__7 
       (.I0(k8[63]),
        .I1(k8[127]),
        .I2(k8[95]),
        .I3(k8[31]),
        .O(\a9/v3 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair250" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[31]_i_1__8 
       (.I0(k9[63]),
        .I1(k9[127]),
        .I2(k9[95]),
        .I3(k9[31]),
        .O(\a10/v3 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair190" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[3]_i_1 
       (.I0(k0[35]),
        .I1(k0[99]),
        .I2(k0[67]),
        .I3(k0[3]),
        .O(\a1/v3 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair161" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[3]_i_1__0 
       (.I0(k1[35]),
        .I1(k1[99]),
        .I2(k1[67]),
        .I3(k1[3]),
        .O(\a2/v3 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair132" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[3]_i_1__1 
       (.I0(k2[35]),
        .I1(k2[99]),
        .I2(k2[67]),
        .I3(k2[3]),
        .O(\a3/v3 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair99" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[3]_i_1__2 
       (.I0(k3[35]),
        .I1(k3[99]),
        .I2(k3[67]),
        .I3(k3[3]),
        .O(\a4/v3 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair70" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[3]_i_1__3 
       (.I0(k4[35]),
        .I1(k4[99]),
        .I2(k4[67]),
        .I3(k4[3]),
        .O(\a5/v3 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair39" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[3]_i_1__4 
       (.I0(k5[35]),
        .I1(k5[99]),
        .I2(k5[67]),
        .I3(k5[3]),
        .O(\a6/v3 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair264" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[3]_i_1__5 
       (.I0(k6[35]),
        .I1(k6[99]),
        .I2(k6[67]),
        .I3(k6[3]),
        .O(\a7/v3 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair313" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[3]_i_1__6 
       (.I0(k7[35]),
        .I1(k7[99]),
        .I2(k7[67]),
        .I3(k7[3]),
        .O(\a8/v3 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair194" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[3]_i_1__7 
       (.I0(k8[35]),
        .I1(k8[99]),
        .I2(k8[67]),
        .I3(k8[3]),
        .O(\a9/v3 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair226" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[3]_i_1__8 
       (.I0(k9[35]),
        .I1(k9[99]),
        .I2(k9[67]),
        .I3(k9[3]),
        .O(\a10/v3 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair189" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[4]_i_1 
       (.I0(k0[36]),
        .I1(k0[100]),
        .I2(k0[68]),
        .I3(k0[4]),
        .O(\a1/v3 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair160" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[4]_i_1__0 
       (.I0(k1[36]),
        .I1(k1[100]),
        .I2(k1[68]),
        .I3(k1[4]),
        .O(\a2/v3 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair131" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[4]_i_1__1 
       (.I0(k2[36]),
        .I1(k2[100]),
        .I2(k2[68]),
        .I3(k2[4]),
        .O(\a3/v3 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair98" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[4]_i_1__2 
       (.I0(k3[36]),
        .I1(k3[100]),
        .I2(k3[68]),
        .I3(k3[4]),
        .O(\a4/v3 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair69" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[4]_i_1__3 
       (.I0(k4[36]),
        .I1(k4[100]),
        .I2(k4[68]),
        .I3(k4[4]),
        .O(\a5/v3 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair40" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[4]_i_1__4 
       (.I0(k5[36]),
        .I1(k5[100]),
        .I2(k5[68]),
        .I3(k5[4]),
        .O(\a6/v3 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair265" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[4]_i_1__5 
       (.I0(k6[36]),
        .I1(k6[100]),
        .I2(k6[68]),
        .I3(k6[4]),
        .O(\a7/v3 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair312" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[4]_i_1__6 
       (.I0(k7[36]),
        .I1(k7[100]),
        .I2(k7[68]),
        .I3(k7[4]),
        .O(\a8/v3 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair195" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[4]_i_1__7 
       (.I0(k8[36]),
        .I1(k8[100]),
        .I2(k8[68]),
        .I3(k8[4]),
        .O(\a9/v3 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair227" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[4]_i_1__8 
       (.I0(k9[36]),
        .I1(k9[100]),
        .I2(k9[68]),
        .I3(k9[4]),
        .O(\a10/v3 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair188" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[5]_i_1 
       (.I0(k0[37]),
        .I1(k0[101]),
        .I2(k0[69]),
        .I3(k0[5]),
        .O(\a1/v3 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair159" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[5]_i_1__0 
       (.I0(k1[37]),
        .I1(k1[101]),
        .I2(k1[69]),
        .I3(k1[5]),
        .O(\a2/v3 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair130" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[5]_i_1__1 
       (.I0(k2[37]),
        .I1(k2[101]),
        .I2(k2[69]),
        .I3(k2[5]),
        .O(\a3/v3 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair97" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[5]_i_1__2 
       (.I0(k3[37]),
        .I1(k3[101]),
        .I2(k3[69]),
        .I3(k3[5]),
        .O(\a4/v3 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair68" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[5]_i_1__3 
       (.I0(k4[37]),
        .I1(k4[101]),
        .I2(k4[69]),
        .I3(k4[5]),
        .O(\a5/v3 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair41" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[5]_i_1__4 
       (.I0(k5[37]),
        .I1(k5[101]),
        .I2(k5[69]),
        .I3(k5[5]),
        .O(\a6/v3 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair266" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[5]_i_1__5 
       (.I0(k6[37]),
        .I1(k6[101]),
        .I2(k6[69]),
        .I3(k6[5]),
        .O(\a7/v3 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair311" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[5]_i_1__6 
       (.I0(k7[37]),
        .I1(k7[101]),
        .I2(k7[69]),
        .I3(k7[5]),
        .O(\a8/v3 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair196" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[5]_i_1__7 
       (.I0(k8[37]),
        .I1(k8[101]),
        .I2(k8[69]),
        .I3(k8[5]),
        .O(\a9/v3 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair228" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[5]_i_1__8 
       (.I0(k9[37]),
        .I1(k9[101]),
        .I2(k9[69]),
        .I3(k9[5]),
        .O(\a10/v3 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair187" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[6]_i_1 
       (.I0(k0[38]),
        .I1(k0[102]),
        .I2(k0[70]),
        .I3(k0[6]),
        .O(\a1/v3 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair158" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[6]_i_1__0 
       (.I0(k1[38]),
        .I1(k1[102]),
        .I2(k1[70]),
        .I3(k1[6]),
        .O(\a2/v3 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair129" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[6]_i_1__1 
       (.I0(k2[38]),
        .I1(k2[102]),
        .I2(k2[70]),
        .I3(k2[6]),
        .O(\a3/v3 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair96" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[6]_i_1__2 
       (.I0(k3[38]),
        .I1(k3[102]),
        .I2(k3[70]),
        .I3(k3[6]),
        .O(\a4/v3 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[6]_i_1__3 
       (.I0(k4[38]),
        .I1(k4[102]),
        .I2(k4[70]),
        .I3(k4[6]),
        .O(\a5/v3 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair42" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[6]_i_1__4 
       (.I0(k5[38]),
        .I1(k5[102]),
        .I2(k5[70]),
        .I3(k5[6]),
        .O(\a6/v3 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair267" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[6]_i_1__5 
       (.I0(k6[38]),
        .I1(k6[102]),
        .I2(k6[70]),
        .I3(k6[6]),
        .O(\a7/v3 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair310" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[6]_i_1__6 
       (.I0(k7[38]),
        .I1(k7[102]),
        .I2(k7[70]),
        .I3(k7[6]),
        .O(\a8/v3 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair197" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[6]_i_1__7 
       (.I0(k8[38]),
        .I1(k8[102]),
        .I2(k8[70]),
        .I3(k8[6]),
        .O(\a9/v3 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair229" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[6]_i_1__8 
       (.I0(k9[38]),
        .I1(k9[102]),
        .I2(k9[70]),
        .I3(k9[6]),
        .O(\a10/v3 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair186" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[7]_i_1 
       (.I0(k0[39]),
        .I1(k0[103]),
        .I2(k0[71]),
        .I3(k0[7]),
        .O(\a1/v3 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair157" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[7]_i_1__0 
       (.I0(k1[39]),
        .I1(k1[103]),
        .I2(k1[71]),
        .I3(k1[7]),
        .O(\a2/v3 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair128" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[7]_i_1__1 
       (.I0(k2[39]),
        .I1(k2[103]),
        .I2(k2[71]),
        .I3(k2[7]),
        .O(\a3/v3 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair95" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[7]_i_1__2 
       (.I0(k3[39]),
        .I1(k3[103]),
        .I2(k3[71]),
        .I3(k3[7]),
        .O(\a4/v3 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair1" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[7]_i_1__3 
       (.I0(k4[39]),
        .I1(k4[103]),
        .I2(k4[71]),
        .I3(k4[7]),
        .O(\a5/v3 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair43" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[7]_i_1__4 
       (.I0(k5[39]),
        .I1(k5[103]),
        .I2(k5[71]),
        .I3(k5[7]),
        .O(\a6/v3 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair268" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[7]_i_1__5 
       (.I0(k6[39]),
        .I1(k6[103]),
        .I2(k6[71]),
        .I3(k6[7]),
        .O(\a7/v3 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair309" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[7]_i_1__6 
       (.I0(k7[39]),
        .I1(k7[103]),
        .I2(k7[71]),
        .I3(k7[7]),
        .O(\a8/v3 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair198" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[7]_i_1__7 
       (.I0(k8[39]),
        .I1(k8[103]),
        .I2(k8[71]),
        .I3(k8[7]),
        .O(\a9/v3 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair230" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[7]_i_1__8 
       (.I0(k9[39]),
        .I1(k9[103]),
        .I2(k9[71]),
        .I3(k9[7]),
        .O(\a10/v3 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair185" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[8]_i_1 
       (.I0(k0[40]),
        .I1(k0[104]),
        .I2(k0[72]),
        .I3(k0[8]),
        .O(\a1/v3 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair156" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[8]_i_1__0 
       (.I0(k1[40]),
        .I1(k1[104]),
        .I2(k1[72]),
        .I3(k1[8]),
        .O(\a2/v3 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair127" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[8]_i_1__1 
       (.I0(k2[40]),
        .I1(k2[104]),
        .I2(k2[72]),
        .I3(k2[8]),
        .O(\a3/v3 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair94" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[8]_i_1__2 
       (.I0(k3[40]),
        .I1(k3[104]),
        .I2(k3[72]),
        .I3(k3[8]),
        .O(\a4/v3 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair0" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[8]_i_1__3 
       (.I0(k4[40]),
        .I1(k4[104]),
        .I2(k4[72]),
        .I3(k4[8]),
        .O(\a5/v3 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair44" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[8]_i_1__4 
       (.I0(k5[40]),
        .I1(k5[104]),
        .I2(k5[72]),
        .I3(k5[8]),
        .O(\a6/v3 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair269" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[8]_i_1__5 
       (.I0(k6[40]),
        .I1(k6[104]),
        .I2(k6[72]),
        .I3(k6[8]),
        .O(\a7/v3 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair308" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[8]_i_1__6 
       (.I0(k7[40]),
        .I1(k7[104]),
        .I2(k7[72]),
        .I3(k7[8]),
        .O(\a8/v3 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair199" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[8]_i_1__7 
       (.I0(k8[40]),
        .I1(k8[104]),
        .I2(k8[72]),
        .I3(k8[8]),
        .O(\a9/v3 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair231" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[8]_i_1__8 
       (.I0(k9[40]),
        .I1(k9[104]),
        .I2(k9[72]),
        .I3(k9[8]),
        .O(\a10/v3 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair184" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[9]_i_1 
       (.I0(k0[41]),
        .I1(k0[105]),
        .I2(k0[73]),
        .I3(k0[9]),
        .O(\a1/v3 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair155" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[9]_i_1__0 
       (.I0(k1[41]),
        .I1(k1[105]),
        .I2(k1[73]),
        .I3(k1[9]),
        .O(\a2/v3 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair126" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[9]_i_1__1 
       (.I0(k2[41]),
        .I1(k2[105]),
        .I2(k2[73]),
        .I3(k2[9]),
        .O(\a3/v3 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair93" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[9]_i_1__2 
       (.I0(k3[41]),
        .I1(k3[105]),
        .I2(k3[73]),
        .I3(k3[9]),
        .O(\a4/v3 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair34" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[9]_i_1__3 
       (.I0(k4[41]),
        .I1(k4[105]),
        .I2(k4[73]),
        .I3(k4[9]),
        .O(\a5/v3 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair45" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[9]_i_1__4 
       (.I0(k5[41]),
        .I1(k5[105]),
        .I2(k5[73]),
        .I3(k5[9]),
        .O(\a6/v3 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair270" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[9]_i_1__5 
       (.I0(k6[41]),
        .I1(k6[105]),
        .I2(k6[73]),
        .I3(k6[9]),
        .O(\a7/v3 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair307" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[9]_i_1__6 
       (.I0(k7[41]),
        .I1(k7[105]),
        .I2(k7[73]),
        .I3(k7[9]),
        .O(\a8/v3 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair200" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[9]_i_1__7 
       (.I0(k8[41]),
        .I1(k8[105]),
        .I2(k8[73]),
        .I3(k8[9]),
        .O(\a9/v3 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair232" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \k3a[9]_i_1__8 
       (.I0(k9[41]),
        .I1(k9[105]),
        .I2(k9[73]),
        .I3(k9[9]),
        .O(\a10/v3 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[0]_i_1 
       (.I0(\a1/k3a [0]),
        .I1(\a1/k4a [0]),
        .O(k0b[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[0]_i_1__0 
       (.I0(\a2/k3a [0]),
        .I1(\a2/k4a [0]),
        .O(k1b[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[0]_i_1__1 
       (.I0(\a3/k3a [0]),
        .I1(\a3/k4a [0]),
        .O(k2b[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[0]_i_1__2 
       (.I0(\a4/k3a [0]),
        .I1(\a4/k4a [0]),
        .O(k3b[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[0]_i_1__3 
       (.I0(\a5/k3a [0]),
        .I1(\a5/k4a [0]),
        .O(k4b[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[0]_i_1__4 
       (.I0(\a6/k3a [0]),
        .I1(\a6/k4a [0]),
        .O(k5b[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[0]_i_1__5 
       (.I0(\a7/k3a [0]),
        .I1(\a7/k4a [0]),
        .O(k6b[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[0]_i_1__6 
       (.I0(\a8/k3a [0]),
        .I1(\a8/k4a [0]),
        .O(k7b[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[0]_i_1__7 
       (.I0(\a9/k3a [0]),
        .I1(\a9/k4a [0]),
        .O(k8b[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[100]_i_1 
       (.I0(\a1/k0a [4]),
        .I1(\a1/k4a [4]),
        .O(k0b[100]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[100]_i_1__0 
       (.I0(\a2/k0a [4]),
        .I1(\a2/k4a [4]),
        .O(k1b[100]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[100]_i_1__1 
       (.I0(\a3/k0a [4]),
        .I1(\a3/k4a [4]),
        .O(k2b[100]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[100]_i_1__2 
       (.I0(\a4/k0a [4]),
        .I1(\a4/k4a [4]),
        .O(k3b[100]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[100]_i_1__3 
       (.I0(\a5/k0a [4]),
        .I1(\a5/k4a [4]),
        .O(k4b[100]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[100]_i_1__4 
       (.I0(\a6/k0a [4]),
        .I1(\a6/k4a [4]),
        .O(k5b[100]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[100]_i_1__5 
       (.I0(\a7/k0a [4]),
        .I1(\a7/k4a [4]),
        .O(k6b[100]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[100]_i_1__6 
       (.I0(\a8/k0a [4]),
        .I1(\a8/k4a [4]),
        .O(k7b[100]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[100]_i_1__7 
       (.I0(\a9/k0a [4]),
        .I1(\a9/k4a [4]),
        .O(k8b[100]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[101]_i_1 
       (.I0(\a1/k0a [5]),
        .I1(\a1/k4a [5]),
        .O(k0b[101]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[101]_i_1__0 
       (.I0(\a2/k0a [5]),
        .I1(\a2/k4a [5]),
        .O(k1b[101]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[101]_i_1__1 
       (.I0(\a3/k0a [5]),
        .I1(\a3/k4a [5]),
        .O(k2b[101]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[101]_i_1__2 
       (.I0(\a4/k0a [5]),
        .I1(\a4/k4a [5]),
        .O(k3b[101]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[101]_i_1__3 
       (.I0(\a5/k0a [5]),
        .I1(\a5/k4a [5]),
        .O(k4b[101]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[101]_i_1__4 
       (.I0(\a6/k0a [5]),
        .I1(\a6/k4a [5]),
        .O(k5b[101]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[101]_i_1__5 
       (.I0(\a7/k0a [5]),
        .I1(\a7/k4a [5]),
        .O(k6b[101]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[101]_i_1__6 
       (.I0(\a8/k0a [5]),
        .I1(\a8/k4a [5]),
        .O(k7b[101]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[101]_i_1__7 
       (.I0(\a9/k0a [5]),
        .I1(\a9/k4a [5]),
        .O(k8b[101]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[102]_i_1 
       (.I0(\a1/k0a [6]),
        .I1(\a1/k4a [6]),
        .O(k0b[102]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[102]_i_1__0 
       (.I0(\a2/k0a [6]),
        .I1(\a2/k4a [6]),
        .O(k1b[102]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[102]_i_1__1 
       (.I0(\a3/k0a [6]),
        .I1(\a3/k4a [6]),
        .O(k2b[102]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[102]_i_1__2 
       (.I0(\a4/k0a [6]),
        .I1(\a4/k4a [6]),
        .O(k3b[102]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[102]_i_1__3 
       (.I0(\a5/k0a [6]),
        .I1(\a5/k4a [6]),
        .O(k4b[102]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[102]_i_1__4 
       (.I0(\a6/k0a [6]),
        .I1(\a6/k4a [6]),
        .O(k5b[102]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[102]_i_1__5 
       (.I0(\a7/k0a [6]),
        .I1(\a7/k4a [6]),
        .O(k6b[102]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[102]_i_1__6 
       (.I0(\a8/k0a [6]),
        .I1(\a8/k4a [6]),
        .O(k7b[102]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[102]_i_1__7 
       (.I0(\a9/k0a [6]),
        .I1(\a9/k4a [6]),
        .O(k8b[102]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[103]_i_1 
       (.I0(\a1/k0a [7]),
        .I1(\a1/k4a [7]),
        .O(k0b[103]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[103]_i_1__0 
       (.I0(\a2/k0a [7]),
        .I1(\a2/k4a [7]),
        .O(k1b[103]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[103]_i_1__1 
       (.I0(\a3/k0a [7]),
        .I1(\a3/k4a [7]),
        .O(k2b[103]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[103]_i_1__2 
       (.I0(\a4/k0a [7]),
        .I1(\a4/k4a [7]),
        .O(k3b[103]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[103]_i_1__3 
       (.I0(\a5/k0a [7]),
        .I1(\a5/k4a [7]),
        .O(k4b[103]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[103]_i_1__4 
       (.I0(\a6/k0a [7]),
        .I1(\a6/k4a [7]),
        .O(k5b[103]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[103]_i_1__5 
       (.I0(\a7/k0a [7]),
        .I1(\a7/k4a [7]),
        .O(k6b[103]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[103]_i_1__6 
       (.I0(\a8/k0a [7]),
        .I1(\a8/k4a [7]),
        .O(k7b[103]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[103]_i_1__7 
       (.I0(\a9/k0a [7]),
        .I1(\a9/k4a [7]),
        .O(k8b[103]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[104]_i_1 
       (.I0(\a1/k0a [8]),
        .I1(\a1/k4a [8]),
        .O(k0b[104]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[104]_i_1__0 
       (.I0(\a2/k0a [8]),
        .I1(\a2/k4a [8]),
        .O(k1b[104]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[104]_i_1__1 
       (.I0(\a3/k0a [8]),
        .I1(\a3/k4a [8]),
        .O(k2b[104]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[104]_i_1__2 
       (.I0(\a4/k0a [8]),
        .I1(\a4/k4a [8]),
        .O(k3b[104]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[104]_i_1__3 
       (.I0(\a5/k0a [8]),
        .I1(\a5/k4a [8]),
        .O(k4b[104]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[104]_i_1__4 
       (.I0(\a6/k0a [8]),
        .I1(\a6/k4a [8]),
        .O(k5b[104]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[104]_i_1__5 
       (.I0(\a7/k0a [8]),
        .I1(\a7/k4a [8]),
        .O(k6b[104]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[104]_i_1__6 
       (.I0(\a8/k0a [8]),
        .I1(\a8/k4a [8]),
        .O(k7b[104]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[104]_i_1__7 
       (.I0(\a9/k0a [8]),
        .I1(\a9/k4a [8]),
        .O(k8b[104]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[105]_i_1 
       (.I0(\a1/k0a [9]),
        .I1(\a1/k4a [9]),
        .O(k0b[105]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[105]_i_1__0 
       (.I0(\a2/k0a [9]),
        .I1(\a2/k4a [9]),
        .O(k1b[105]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[105]_i_1__1 
       (.I0(\a3/k0a [9]),
        .I1(\a3/k4a [9]),
        .O(k2b[105]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[105]_i_1__2 
       (.I0(\a4/k0a [9]),
        .I1(\a4/k4a [9]),
        .O(k3b[105]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[105]_i_1__3 
       (.I0(\a5/k0a [9]),
        .I1(\a5/k4a [9]),
        .O(k4b[105]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[105]_i_1__4 
       (.I0(\a6/k0a [9]),
        .I1(\a6/k4a [9]),
        .O(k5b[105]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[105]_i_1__5 
       (.I0(\a7/k0a [9]),
        .I1(\a7/k4a [9]),
        .O(k6b[105]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[105]_i_1__6 
       (.I0(\a8/k0a [9]),
        .I1(\a8/k4a [9]),
        .O(k7b[105]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[105]_i_1__7 
       (.I0(\a9/k0a [9]),
        .I1(\a9/k4a [9]),
        .O(k8b[105]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[106]_i_1 
       (.I0(\a1/k0a [10]),
        .I1(\a1/k4a [10]),
        .O(k0b[106]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[106]_i_1__0 
       (.I0(\a2/k0a [10]),
        .I1(\a2/k4a [10]),
        .O(k1b[106]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[106]_i_1__1 
       (.I0(\a3/k0a [10]),
        .I1(\a3/k4a [10]),
        .O(k2b[106]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[106]_i_1__2 
       (.I0(\a4/k0a [10]),
        .I1(\a4/k4a [10]),
        .O(k3b[106]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[106]_i_1__3 
       (.I0(\a5/k0a [10]),
        .I1(\a5/k4a [10]),
        .O(k4b[106]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[106]_i_1__4 
       (.I0(\a6/k0a [10]),
        .I1(\a6/k4a [10]),
        .O(k5b[106]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[106]_i_1__5 
       (.I0(\a7/k0a [10]),
        .I1(\a7/k4a [10]),
        .O(k6b[106]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[106]_i_1__6 
       (.I0(\a8/k0a [10]),
        .I1(\a8/k4a [10]),
        .O(k7b[106]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[106]_i_1__7 
       (.I0(\a9/k0a [10]),
        .I1(\a9/k4a [10]),
        .O(k8b[106]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[107]_i_1 
       (.I0(\a1/k0a [11]),
        .I1(\a1/k4a [11]),
        .O(k0b[107]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[107]_i_1__0 
       (.I0(\a2/k0a [11]),
        .I1(\a2/k4a [11]),
        .O(k1b[107]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[107]_i_1__1 
       (.I0(\a3/k0a [11]),
        .I1(\a3/k4a [11]),
        .O(k2b[107]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[107]_i_1__2 
       (.I0(\a4/k0a [11]),
        .I1(\a4/k4a [11]),
        .O(k3b[107]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[107]_i_1__3 
       (.I0(\a5/k0a [11]),
        .I1(\a5/k4a [11]),
        .O(k4b[107]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[107]_i_1__4 
       (.I0(\a6/k0a [11]),
        .I1(\a6/k4a [11]),
        .O(k5b[107]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[107]_i_1__5 
       (.I0(\a7/k0a [11]),
        .I1(\a7/k4a [11]),
        .O(k6b[107]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[107]_i_1__6 
       (.I0(\a8/k0a [11]),
        .I1(\a8/k4a [11]),
        .O(k7b[107]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[107]_i_1__7 
       (.I0(\a9/k0a [11]),
        .I1(\a9/k4a [11]),
        .O(k8b[107]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[108]_i_1 
       (.I0(\a1/k0a [12]),
        .I1(\a1/k4a [12]),
        .O(k0b[108]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[108]_i_1__0 
       (.I0(\a2/k0a [12]),
        .I1(\a2/k4a [12]),
        .O(k1b[108]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[108]_i_1__1 
       (.I0(\a3/k0a [12]),
        .I1(\a3/k4a [12]),
        .O(k2b[108]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[108]_i_1__2 
       (.I0(\a4/k0a [12]),
        .I1(\a4/k4a [12]),
        .O(k3b[108]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[108]_i_1__3 
       (.I0(\a5/k0a [12]),
        .I1(\a5/k4a [12]),
        .O(k4b[108]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[108]_i_1__4 
       (.I0(\a6/k0a [12]),
        .I1(\a6/k4a [12]),
        .O(k5b[108]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[108]_i_1__5 
       (.I0(\a7/k0a [12]),
        .I1(\a7/k4a [12]),
        .O(k6b[108]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[108]_i_1__6 
       (.I0(\a8/k0a [12]),
        .I1(\a8/k4a [12]),
        .O(k7b[108]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[108]_i_1__7 
       (.I0(\a9/k0a [12]),
        .I1(\a9/k4a [12]),
        .O(k8b[108]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[109]_i_1 
       (.I0(\a1/k0a [13]),
        .I1(\a1/k4a [13]),
        .O(k0b[109]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[109]_i_1__0 
       (.I0(\a2/k0a [13]),
        .I1(\a2/k4a [13]),
        .O(k1b[109]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[109]_i_1__1 
       (.I0(\a3/k0a [13]),
        .I1(\a3/k4a [13]),
        .O(k2b[109]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[109]_i_1__2 
       (.I0(\a4/k0a [13]),
        .I1(\a4/k4a [13]),
        .O(k3b[109]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[109]_i_1__3 
       (.I0(\a5/k0a [13]),
        .I1(\a5/k4a [13]),
        .O(k4b[109]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[109]_i_1__4 
       (.I0(\a6/k0a [13]),
        .I1(\a6/k4a [13]),
        .O(k5b[109]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[109]_i_1__5 
       (.I0(\a7/k0a [13]),
        .I1(\a7/k4a [13]),
        .O(k6b[109]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[109]_i_1__6 
       (.I0(\a8/k0a [13]),
        .I1(\a8/k4a [13]),
        .O(k7b[109]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[109]_i_1__7 
       (.I0(\a9/k0a [13]),
        .I1(\a9/k4a [13]),
        .O(k8b[109]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[10]_i_1 
       (.I0(\a1/k3a [10]),
        .I1(\a1/k4a [10]),
        .O(k0b[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[10]_i_1__0 
       (.I0(\a2/k3a [10]),
        .I1(\a2/k4a [10]),
        .O(k1b[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[10]_i_1__1 
       (.I0(\a3/k3a [10]),
        .I1(\a3/k4a [10]),
        .O(k2b[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[10]_i_1__2 
       (.I0(\a4/k3a [10]),
        .I1(\a4/k4a [10]),
        .O(k3b[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[10]_i_1__3 
       (.I0(\a5/k3a [10]),
        .I1(\a5/k4a [10]),
        .O(k4b[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[10]_i_1__4 
       (.I0(\a6/k3a [10]),
        .I1(\a6/k4a [10]),
        .O(k5b[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[10]_i_1__5 
       (.I0(\a7/k3a [10]),
        .I1(\a7/k4a [10]),
        .O(k6b[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[10]_i_1__6 
       (.I0(\a8/k3a [10]),
        .I1(\a8/k4a [10]),
        .O(k7b[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[10]_i_1__7 
       (.I0(\a9/k3a [10]),
        .I1(\a9/k4a [10]),
        .O(k8b[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[110]_i_1 
       (.I0(\a1/k0a [14]),
        .I1(\a1/k4a [14]),
        .O(k0b[110]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[110]_i_1__0 
       (.I0(\a2/k0a [14]),
        .I1(\a2/k4a [14]),
        .O(k1b[110]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[110]_i_1__1 
       (.I0(\a3/k0a [14]),
        .I1(\a3/k4a [14]),
        .O(k2b[110]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[110]_i_1__2 
       (.I0(\a4/k0a [14]),
        .I1(\a4/k4a [14]),
        .O(k3b[110]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[110]_i_1__3 
       (.I0(\a5/k0a [14]),
        .I1(\a5/k4a [14]),
        .O(k4b[110]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[110]_i_1__4 
       (.I0(\a6/k0a [14]),
        .I1(\a6/k4a [14]),
        .O(k5b[110]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[110]_i_1__5 
       (.I0(\a7/k0a [14]),
        .I1(\a7/k4a [14]),
        .O(k6b[110]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[110]_i_1__6 
       (.I0(\a8/k0a [14]),
        .I1(\a8/k4a [14]),
        .O(k7b[110]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[110]_i_1__7 
       (.I0(\a9/k0a [14]),
        .I1(\a9/k4a [14]),
        .O(k8b[110]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[111]_i_1 
       (.I0(\a1/k0a [15]),
        .I1(\a1/k4a [15]),
        .O(k0b[111]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[111]_i_1__0 
       (.I0(\a2/k0a [15]),
        .I1(\a2/k4a [15]),
        .O(k1b[111]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[111]_i_1__1 
       (.I0(\a3/k0a [15]),
        .I1(\a3/k4a [15]),
        .O(k2b[111]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[111]_i_1__2 
       (.I0(\a4/k0a [15]),
        .I1(\a4/k4a [15]),
        .O(k3b[111]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[111]_i_1__3 
       (.I0(\a5/k0a [15]),
        .I1(\a5/k4a [15]),
        .O(k4b[111]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[111]_i_1__4 
       (.I0(\a6/k0a [15]),
        .I1(\a6/k4a [15]),
        .O(k5b[111]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[111]_i_1__5 
       (.I0(\a7/k0a [15]),
        .I1(\a7/k4a [15]),
        .O(k6b[111]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[111]_i_1__6 
       (.I0(\a8/k0a [15]),
        .I1(\a8/k4a [15]),
        .O(k7b[111]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[111]_i_1__7 
       (.I0(\a9/k0a [15]),
        .I1(\a9/k4a [15]),
        .O(k8b[111]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[112]_i_1 
       (.I0(\a1/k0a [16]),
        .I1(\a1/k4a [16]),
        .O(k0b[112]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[112]_i_1__0 
       (.I0(\a2/k0a [16]),
        .I1(\a2/k4a [16]),
        .O(k1b[112]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[112]_i_1__1 
       (.I0(\a3/k0a [16]),
        .I1(\a3/k4a [16]),
        .O(k2b[112]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[112]_i_1__2 
       (.I0(\a4/k0a [16]),
        .I1(\a4/k4a [16]),
        .O(k3b[112]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[112]_i_1__3 
       (.I0(\a5/k0a [16]),
        .I1(\a5/k4a [16]),
        .O(k4b[112]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[112]_i_1__4 
       (.I0(\a6/k0a [16]),
        .I1(\a6/k4a [16]),
        .O(k5b[112]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[112]_i_1__5 
       (.I0(\a7/k0a [16]),
        .I1(\a7/k4a [16]),
        .O(k6b[112]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[112]_i_1__6 
       (.I0(\a8/k0a [16]),
        .I1(\a8/k4a [16]),
        .O(k7b[112]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[112]_i_1__7 
       (.I0(\a9/k0a [16]),
        .I1(\a9/k4a [16]),
        .O(k8b[112]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[113]_i_1 
       (.I0(\a1/k0a [17]),
        .I1(\a1/k4a [17]),
        .O(k0b[113]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[113]_i_1__0 
       (.I0(\a2/k0a [17]),
        .I1(\a2/k4a [17]),
        .O(k1b[113]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[113]_i_1__1 
       (.I0(\a3/k0a [17]),
        .I1(\a3/k4a [17]),
        .O(k2b[113]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[113]_i_1__2 
       (.I0(\a4/k0a [17]),
        .I1(\a4/k4a [17]),
        .O(k3b[113]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[113]_i_1__3 
       (.I0(\a5/k0a [17]),
        .I1(\a5/k4a [17]),
        .O(k4b[113]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[113]_i_1__4 
       (.I0(\a6/k0a [17]),
        .I1(\a6/k4a [17]),
        .O(k5b[113]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[113]_i_1__5 
       (.I0(\a7/k0a [17]),
        .I1(\a7/k4a [17]),
        .O(k6b[113]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[113]_i_1__6 
       (.I0(\a8/k0a [17]),
        .I1(\a8/k4a [17]),
        .O(k7b[113]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[113]_i_1__7 
       (.I0(\a9/k0a [17]),
        .I1(\a9/k4a [17]),
        .O(k8b[113]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[114]_i_1 
       (.I0(\a1/k0a [18]),
        .I1(\a1/k4a [18]),
        .O(k0b[114]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[114]_i_1__0 
       (.I0(\a2/k0a [18]),
        .I1(\a2/k4a [18]),
        .O(k1b[114]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[114]_i_1__1 
       (.I0(\a3/k0a [18]),
        .I1(\a3/k4a [18]),
        .O(k2b[114]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[114]_i_1__2 
       (.I0(\a4/k0a [18]),
        .I1(\a4/k4a [18]),
        .O(k3b[114]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[114]_i_1__3 
       (.I0(\a5/k0a [18]),
        .I1(\a5/k4a [18]),
        .O(k4b[114]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[114]_i_1__4 
       (.I0(\a6/k0a [18]),
        .I1(\a6/k4a [18]),
        .O(k5b[114]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[114]_i_1__5 
       (.I0(\a7/k0a [18]),
        .I1(\a7/k4a [18]),
        .O(k6b[114]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[114]_i_1__6 
       (.I0(\a8/k0a [18]),
        .I1(\a8/k4a [18]),
        .O(k7b[114]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[114]_i_1__7 
       (.I0(\a9/k0a [18]),
        .I1(\a9/k4a [18]),
        .O(k8b[114]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[115]_i_1 
       (.I0(\a1/k0a [19]),
        .I1(\a1/k4a [19]),
        .O(k0b[115]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[115]_i_1__0 
       (.I0(\a2/k0a [19]),
        .I1(\a2/k4a [19]),
        .O(k1b[115]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[115]_i_1__1 
       (.I0(\a3/k0a [19]),
        .I1(\a3/k4a [19]),
        .O(k2b[115]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[115]_i_1__2 
       (.I0(\a4/k0a [19]),
        .I1(\a4/k4a [19]),
        .O(k3b[115]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[115]_i_1__3 
       (.I0(\a5/k0a [19]),
        .I1(\a5/k4a [19]),
        .O(k4b[115]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[115]_i_1__4 
       (.I0(\a6/k0a [19]),
        .I1(\a6/k4a [19]),
        .O(k5b[115]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[115]_i_1__5 
       (.I0(\a7/k0a [19]),
        .I1(\a7/k4a [19]),
        .O(k6b[115]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[115]_i_1__6 
       (.I0(\a8/k0a [19]),
        .I1(\a8/k4a [19]),
        .O(k7b[115]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[115]_i_1__7 
       (.I0(\a9/k0a [19]),
        .I1(\a9/k4a [19]),
        .O(k8b[115]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[116]_i_1 
       (.I0(\a1/k0a [20]),
        .I1(\a1/k4a [20]),
        .O(k0b[116]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[116]_i_1__0 
       (.I0(\a2/k0a [20]),
        .I1(\a2/k4a [20]),
        .O(k1b[116]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[116]_i_1__1 
       (.I0(\a3/k0a [20]),
        .I1(\a3/k4a [20]),
        .O(k2b[116]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[116]_i_1__2 
       (.I0(\a4/k0a [20]),
        .I1(\a4/k4a [20]),
        .O(k3b[116]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[116]_i_1__3 
       (.I0(\a5/k0a [20]),
        .I1(\a5/k4a [20]),
        .O(k4b[116]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[116]_i_1__4 
       (.I0(\a6/k0a [20]),
        .I1(\a6/k4a [20]),
        .O(k5b[116]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[116]_i_1__5 
       (.I0(\a7/k0a [20]),
        .I1(\a7/k4a [20]),
        .O(k6b[116]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[116]_i_1__6 
       (.I0(\a8/k0a [20]),
        .I1(\a8/k4a [20]),
        .O(k7b[116]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[116]_i_1__7 
       (.I0(\a9/k0a [20]),
        .I1(\a9/k4a [20]),
        .O(k8b[116]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[117]_i_1 
       (.I0(\a1/k0a [21]),
        .I1(\a1/k4a [21]),
        .O(k0b[117]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[117]_i_1__0 
       (.I0(\a2/k0a [21]),
        .I1(\a2/k4a [21]),
        .O(k1b[117]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[117]_i_1__1 
       (.I0(\a3/k0a [21]),
        .I1(\a3/k4a [21]),
        .O(k2b[117]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[117]_i_1__2 
       (.I0(\a4/k0a [21]),
        .I1(\a4/k4a [21]),
        .O(k3b[117]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[117]_i_1__3 
       (.I0(\a5/k0a [21]),
        .I1(\a5/k4a [21]),
        .O(k4b[117]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[117]_i_1__4 
       (.I0(\a6/k0a [21]),
        .I1(\a6/k4a [21]),
        .O(k5b[117]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[117]_i_1__5 
       (.I0(\a7/k0a [21]),
        .I1(\a7/k4a [21]),
        .O(k6b[117]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[117]_i_1__6 
       (.I0(\a8/k0a [21]),
        .I1(\a8/k4a [21]),
        .O(k7b[117]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[117]_i_1__7 
       (.I0(\a9/k0a [21]),
        .I1(\a9/k4a [21]),
        .O(k8b[117]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[118]_i_1 
       (.I0(\a1/k0a [22]),
        .I1(\a1/k4a [22]),
        .O(k0b[118]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[118]_i_1__0 
       (.I0(\a2/k0a [22]),
        .I1(\a2/k4a [22]),
        .O(k1b[118]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[118]_i_1__1 
       (.I0(\a3/k0a [22]),
        .I1(\a3/k4a [22]),
        .O(k2b[118]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[118]_i_1__2 
       (.I0(\a4/k0a [22]),
        .I1(\a4/k4a [22]),
        .O(k3b[118]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[118]_i_1__3 
       (.I0(\a5/k0a [22]),
        .I1(\a5/k4a [22]),
        .O(k4b[118]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[118]_i_1__4 
       (.I0(\a6/k0a [22]),
        .I1(\a6/k4a [22]),
        .O(k5b[118]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[118]_i_1__5 
       (.I0(\a7/k0a [22]),
        .I1(\a7/k4a [22]),
        .O(k6b[118]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[118]_i_1__6 
       (.I0(\a8/k0a [22]),
        .I1(\a8/k4a [22]),
        .O(k7b[118]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[118]_i_1__7 
       (.I0(\a9/k0a [22]),
        .I1(\a9/k4a [22]),
        .O(k8b[118]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[119]_i_1 
       (.I0(\a1/k0a [23]),
        .I1(\a1/k4a [23]),
        .O(k0b[119]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[119]_i_1__0 
       (.I0(\a2/k0a [23]),
        .I1(\a2/k4a [23]),
        .O(k1b[119]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[119]_i_1__1 
       (.I0(\a3/k0a [23]),
        .I1(\a3/k4a [23]),
        .O(k2b[119]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[119]_i_1__2 
       (.I0(\a4/k0a [23]),
        .I1(\a4/k4a [23]),
        .O(k3b[119]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[119]_i_1__3 
       (.I0(\a5/k0a [23]),
        .I1(\a5/k4a [23]),
        .O(k4b[119]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[119]_i_1__4 
       (.I0(\a6/k0a [23]),
        .I1(\a6/k4a [23]),
        .O(k5b[119]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[119]_i_1__5 
       (.I0(\a7/k0a [23]),
        .I1(\a7/k4a [23]),
        .O(k6b[119]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[119]_i_1__6 
       (.I0(\a8/k0a [23]),
        .I1(\a8/k4a [23]),
        .O(k7b[119]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[119]_i_1__7 
       (.I0(\a9/k0a [23]),
        .I1(\a9/k4a [23]),
        .O(k8b[119]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[11]_i_1 
       (.I0(\a1/k3a [11]),
        .I1(\a1/k4a [11]),
        .O(k0b[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[11]_i_1__0 
       (.I0(\a2/k3a [11]),
        .I1(\a2/k4a [11]),
        .O(k1b[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[11]_i_1__1 
       (.I0(\a3/k3a [11]),
        .I1(\a3/k4a [11]),
        .O(k2b[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[11]_i_1__2 
       (.I0(\a4/k3a [11]),
        .I1(\a4/k4a [11]),
        .O(k3b[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[11]_i_1__3 
       (.I0(\a5/k3a [11]),
        .I1(\a5/k4a [11]),
        .O(k4b[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[11]_i_1__4 
       (.I0(\a6/k3a [11]),
        .I1(\a6/k4a [11]),
        .O(k5b[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[11]_i_1__5 
       (.I0(\a7/k3a [11]),
        .I1(\a7/k4a [11]),
        .O(k6b[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[11]_i_1__6 
       (.I0(\a8/k3a [11]),
        .I1(\a8/k4a [11]),
        .O(k7b[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[11]_i_1__7 
       (.I0(\a9/k3a [11]),
        .I1(\a9/k4a [11]),
        .O(k8b[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[120]_i_1 
       (.I0(\a1/k0a [24]),
        .I1(\a1/k4a [24]),
        .O(k0b[120]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[120]_i_1__0 
       (.I0(\a2/k0a [24]),
        .I1(\a2/k4a [24]),
        .O(k1b[120]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[120]_i_1__1 
       (.I0(\a3/k0a [24]),
        .I1(\a3/k4a [24]),
        .O(k2b[120]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[120]_i_1__2 
       (.I0(\a4/k0a [24]),
        .I1(\a4/k4a [24]),
        .O(k3b[120]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[120]_i_1__3 
       (.I0(\a5/k0a [24]),
        .I1(\a5/k4a [24]),
        .O(k4b[120]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[120]_i_1__4 
       (.I0(\a6/k0a [24]),
        .I1(\a6/k4a [24]),
        .O(k5b[120]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[120]_i_1__5 
       (.I0(\a7/k0a [24]),
        .I1(\a7/k4a [24]),
        .O(k6b[120]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[120]_i_1__6 
       (.I0(\a8/k0a [24]),
        .I1(\a8/k4a [24]),
        .O(k7b[120]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[120]_i_1__7 
       (.I0(\a9/k0a [24]),
        .I1(\a9/k4a [24]),
        .O(k8b[120]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[121]_i_1 
       (.I0(\a1/k0a [25]),
        .I1(\a1/k4a [25]),
        .O(k0b[121]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[121]_i_1__0 
       (.I0(\a2/k0a [25]),
        .I1(\a2/k4a [25]),
        .O(k1b[121]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[121]_i_1__1 
       (.I0(\a3/k0a [25]),
        .I1(\a3/k4a [25]),
        .O(k2b[121]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[121]_i_1__2 
       (.I0(\a4/k0a [25]),
        .I1(\a4/k4a [25]),
        .O(k3b[121]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[121]_i_1__3 
       (.I0(\a5/k0a [25]),
        .I1(\a5/k4a [25]),
        .O(k4b[121]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[121]_i_1__4 
       (.I0(\a6/k0a [25]),
        .I1(\a6/k4a [25]),
        .O(k5b[121]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[121]_i_1__5 
       (.I0(\a7/k0a [25]),
        .I1(\a7/k4a [25]),
        .O(k6b[121]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[121]_i_1__6 
       (.I0(\a8/k0a [25]),
        .I1(\a8/k4a [25]),
        .O(k7b[121]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[121]_i_1__7 
       (.I0(\a9/k0a [25]),
        .I1(\a9/k4a [25]),
        .O(k8b[121]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[122]_i_1 
       (.I0(\a1/k0a [26]),
        .I1(\a1/k4a [26]),
        .O(k0b[122]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[122]_i_1__0 
       (.I0(\a2/k0a [26]),
        .I1(\a2/k4a [26]),
        .O(k1b[122]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[122]_i_1__1 
       (.I0(\a3/k0a [26]),
        .I1(\a3/k4a [26]),
        .O(k2b[122]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[122]_i_1__2 
       (.I0(\a4/k0a [26]),
        .I1(\a4/k4a [26]),
        .O(k3b[122]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[122]_i_1__3 
       (.I0(\a5/k0a [26]),
        .I1(\a5/k4a [26]),
        .O(k4b[122]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[122]_i_1__4 
       (.I0(\a6/k0a [26]),
        .I1(\a6/k4a [26]),
        .O(k5b[122]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[122]_i_1__5 
       (.I0(\a7/k0a [26]),
        .I1(\a7/k4a [26]),
        .O(k6b[122]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[122]_i_1__6 
       (.I0(\a8/k0a [26]),
        .I1(\a8/k4a [26]),
        .O(k7b[122]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[122]_i_1__7 
       (.I0(\a9/k0a [26]),
        .I1(\a9/k4a [26]),
        .O(k8b[122]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[123]_i_1 
       (.I0(\a1/k0a [27]),
        .I1(\a1/k4a [27]),
        .O(k0b[123]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[123]_i_1__0 
       (.I0(\a2/k0a [27]),
        .I1(\a2/k4a [27]),
        .O(k1b[123]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[123]_i_1__1 
       (.I0(\a3/k0a [27]),
        .I1(\a3/k4a [27]),
        .O(k2b[123]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[123]_i_1__2 
       (.I0(\a4/k0a [27]),
        .I1(\a4/k4a [27]),
        .O(k3b[123]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[123]_i_1__3 
       (.I0(\a5/k0a [27]),
        .I1(\a5/k4a [27]),
        .O(k4b[123]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[123]_i_1__4 
       (.I0(\a6/k0a [27]),
        .I1(\a6/k4a [27]),
        .O(k5b[123]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[123]_i_1__5 
       (.I0(\a7/k0a [27]),
        .I1(\a7/k4a [27]),
        .O(k6b[123]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[123]_i_1__6 
       (.I0(\a8/k0a [27]),
        .I1(\a8/k4a [27]),
        .O(k7b[123]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[123]_i_1__7 
       (.I0(\a9/k0a [27]),
        .I1(\a9/k4a [27]),
        .O(k8b[123]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[124]_i_1 
       (.I0(\a1/k0a [28]),
        .I1(\a1/k4a [28]),
        .O(k0b[124]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[124]_i_1__0 
       (.I0(\a2/k0a [28]),
        .I1(\a2/k4a [28]),
        .O(k1b[124]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[124]_i_1__1 
       (.I0(\a3/k0a [28]),
        .I1(\a3/k4a [28]),
        .O(k2b[124]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[124]_i_1__2 
       (.I0(\a4/k0a [28]),
        .I1(\a4/k4a [28]),
        .O(k3b[124]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[124]_i_1__3 
       (.I0(\a5/k0a [28]),
        .I1(\a5/k4a [28]),
        .O(k4b[124]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[124]_i_1__4 
       (.I0(\a6/k0a [28]),
        .I1(\a6/k4a [28]),
        .O(k5b[124]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[124]_i_1__5 
       (.I0(\a7/k0a [28]),
        .I1(\a7/k4a [28]),
        .O(k6b[124]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[124]_i_1__6 
       (.I0(\a8/k0a [28]),
        .I1(\a8/k4a [28]),
        .O(k7b[124]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[124]_i_1__7 
       (.I0(\a9/k0a [28]),
        .I1(\a9/k4a [28]),
        .O(k8b[124]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[125]_i_1 
       (.I0(\a1/k0a [29]),
        .I1(\a1/k4a [29]),
        .O(k0b[125]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[125]_i_1__0 
       (.I0(\a2/k0a [29]),
        .I1(\a2/k4a [29]),
        .O(k1b[125]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[125]_i_1__1 
       (.I0(\a3/k0a [29]),
        .I1(\a3/k4a [29]),
        .O(k2b[125]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[125]_i_1__2 
       (.I0(\a4/k0a [29]),
        .I1(\a4/k4a [29]),
        .O(k3b[125]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[125]_i_1__3 
       (.I0(\a5/k0a [29]),
        .I1(\a5/k4a [29]),
        .O(k4b[125]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[125]_i_1__4 
       (.I0(\a6/k0a [29]),
        .I1(\a6/k4a [29]),
        .O(k5b[125]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[125]_i_1__5 
       (.I0(\a7/k0a [29]),
        .I1(\a7/k4a [29]),
        .O(k6b[125]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[125]_i_1__6 
       (.I0(\a8/k0a [29]),
        .I1(\a8/k4a [29]),
        .O(k7b[125]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[125]_i_1__7 
       (.I0(\a9/k0a [29]),
        .I1(\a9/k4a [29]),
        .O(k8b[125]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[126]_i_1 
       (.I0(\a1/k0a [30]),
        .I1(\a1/k4a [30]),
        .O(k0b[126]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[126]_i_1__0 
       (.I0(\a2/k0a [30]),
        .I1(\a2/k4a [30]),
        .O(k1b[126]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[126]_i_1__1 
       (.I0(\a3/k0a [30]),
        .I1(\a3/k4a [30]),
        .O(k2b[126]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[126]_i_1__2 
       (.I0(\a4/k0a [30]),
        .I1(\a4/k4a [30]),
        .O(k3b[126]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[126]_i_1__3 
       (.I0(\a5/k0a [30]),
        .I1(\a5/k4a [30]),
        .O(k4b[126]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[126]_i_1__4 
       (.I0(\a6/k0a [30]),
        .I1(\a6/k4a [30]),
        .O(k5b[126]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[126]_i_1__5 
       (.I0(\a7/k0a [30]),
        .I1(\a7/k4a [30]),
        .O(k6b[126]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[126]_i_1__6 
       (.I0(\a8/k0a [30]),
        .I1(\a8/k4a [30]),
        .O(k7b[126]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[126]_i_1__7 
       (.I0(\a9/k0a [30]),
        .I1(\a9/k4a [30]),
        .O(k8b[126]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[127]_i_1 
       (.I0(\a1/k0a [31]),
        .I1(\a1/k4a [31]),
        .O(k0b[127]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[127]_i_1__0 
       (.I0(\a2/k0a [31]),
        .I1(\a2/k4a [31]),
        .O(k1b[127]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[127]_i_1__1 
       (.I0(\a3/k0a [31]),
        .I1(\a3/k4a [31]),
        .O(k2b[127]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[127]_i_1__2 
       (.I0(\a4/k0a [31]),
        .I1(\a4/k4a [31]),
        .O(k3b[127]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[127]_i_1__3 
       (.I0(\a5/k0a [31]),
        .I1(\a5/k4a [31]),
        .O(k4b[127]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[127]_i_1__4 
       (.I0(\a6/k0a [31]),
        .I1(\a6/k4a [31]),
        .O(k5b[127]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[127]_i_1__5 
       (.I0(\a7/k0a [31]),
        .I1(\a7/k4a [31]),
        .O(k6b[127]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[127]_i_1__6 
       (.I0(\a8/k0a [31]),
        .I1(\a8/k4a [31]),
        .O(k7b[127]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[127]_i_1__7 
       (.I0(\a9/k0a [31]),
        .I1(\a9/k4a [31]),
        .O(k8b[127]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[12]_i_1 
       (.I0(\a1/k3a [12]),
        .I1(\a1/k4a [12]),
        .O(k0b[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[12]_i_1__0 
       (.I0(\a2/k3a [12]),
        .I1(\a2/k4a [12]),
        .O(k1b[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[12]_i_1__1 
       (.I0(\a3/k3a [12]),
        .I1(\a3/k4a [12]),
        .O(k2b[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[12]_i_1__2 
       (.I0(\a4/k3a [12]),
        .I1(\a4/k4a [12]),
        .O(k3b[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[12]_i_1__3 
       (.I0(\a5/k3a [12]),
        .I1(\a5/k4a [12]),
        .O(k4b[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[12]_i_1__4 
       (.I0(\a6/k3a [12]),
        .I1(\a6/k4a [12]),
        .O(k5b[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[12]_i_1__5 
       (.I0(\a7/k3a [12]),
        .I1(\a7/k4a [12]),
        .O(k6b[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[12]_i_1__6 
       (.I0(\a8/k3a [12]),
        .I1(\a8/k4a [12]),
        .O(k7b[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[12]_i_1__7 
       (.I0(\a9/k3a [12]),
        .I1(\a9/k4a [12]),
        .O(k8b[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[13]_i_1 
       (.I0(\a1/k3a [13]),
        .I1(\a1/k4a [13]),
        .O(k0b[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[13]_i_1__0 
       (.I0(\a2/k3a [13]),
        .I1(\a2/k4a [13]),
        .O(k1b[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[13]_i_1__1 
       (.I0(\a3/k3a [13]),
        .I1(\a3/k4a [13]),
        .O(k2b[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[13]_i_1__2 
       (.I0(\a4/k3a [13]),
        .I1(\a4/k4a [13]),
        .O(k3b[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[13]_i_1__3 
       (.I0(\a5/k3a [13]),
        .I1(\a5/k4a [13]),
        .O(k4b[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[13]_i_1__4 
       (.I0(\a6/k3a [13]),
        .I1(\a6/k4a [13]),
        .O(k5b[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[13]_i_1__5 
       (.I0(\a7/k3a [13]),
        .I1(\a7/k4a [13]),
        .O(k6b[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[13]_i_1__6 
       (.I0(\a8/k3a [13]),
        .I1(\a8/k4a [13]),
        .O(k7b[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[13]_i_1__7 
       (.I0(\a9/k3a [13]),
        .I1(\a9/k4a [13]),
        .O(k8b[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[14]_i_1 
       (.I0(\a1/k3a [14]),
        .I1(\a1/k4a [14]),
        .O(k0b[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[14]_i_1__0 
       (.I0(\a2/k3a [14]),
        .I1(\a2/k4a [14]),
        .O(k1b[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[14]_i_1__1 
       (.I0(\a3/k3a [14]),
        .I1(\a3/k4a [14]),
        .O(k2b[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[14]_i_1__2 
       (.I0(\a4/k3a [14]),
        .I1(\a4/k4a [14]),
        .O(k3b[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[14]_i_1__3 
       (.I0(\a5/k3a [14]),
        .I1(\a5/k4a [14]),
        .O(k4b[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[14]_i_1__4 
       (.I0(\a6/k3a [14]),
        .I1(\a6/k4a [14]),
        .O(k5b[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[14]_i_1__5 
       (.I0(\a7/k3a [14]),
        .I1(\a7/k4a [14]),
        .O(k6b[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[14]_i_1__6 
       (.I0(\a8/k3a [14]),
        .I1(\a8/k4a [14]),
        .O(k7b[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[14]_i_1__7 
       (.I0(\a9/k3a [14]),
        .I1(\a9/k4a [14]),
        .O(k8b[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[15]_i_1 
       (.I0(\a1/k3a [15]),
        .I1(\a1/k4a [15]),
        .O(k0b[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[15]_i_1__0 
       (.I0(\a2/k3a [15]),
        .I1(\a2/k4a [15]),
        .O(k1b[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[15]_i_1__1 
       (.I0(\a3/k3a [15]),
        .I1(\a3/k4a [15]),
        .O(k2b[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[15]_i_1__2 
       (.I0(\a4/k3a [15]),
        .I1(\a4/k4a [15]),
        .O(k3b[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[15]_i_1__3 
       (.I0(\a5/k3a [15]),
        .I1(\a5/k4a [15]),
        .O(k4b[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[15]_i_1__4 
       (.I0(\a6/k3a [15]),
        .I1(\a6/k4a [15]),
        .O(k5b[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[15]_i_1__5 
       (.I0(\a7/k3a [15]),
        .I1(\a7/k4a [15]),
        .O(k6b[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[15]_i_1__6 
       (.I0(\a8/k3a [15]),
        .I1(\a8/k4a [15]),
        .O(k7b[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[15]_i_1__7 
       (.I0(\a9/k3a [15]),
        .I1(\a9/k4a [15]),
        .O(k8b[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[16]_i_1 
       (.I0(\a1/k3a [16]),
        .I1(\a1/k4a [16]),
        .O(k0b[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[16]_i_1__0 
       (.I0(\a2/k3a [16]),
        .I1(\a2/k4a [16]),
        .O(k1b[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[16]_i_1__1 
       (.I0(\a3/k3a [16]),
        .I1(\a3/k4a [16]),
        .O(k2b[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[16]_i_1__2 
       (.I0(\a4/k3a [16]),
        .I1(\a4/k4a [16]),
        .O(k3b[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[16]_i_1__3 
       (.I0(\a5/k3a [16]),
        .I1(\a5/k4a [16]),
        .O(k4b[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[16]_i_1__4 
       (.I0(\a6/k3a [16]),
        .I1(\a6/k4a [16]),
        .O(k5b[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[16]_i_1__5 
       (.I0(\a7/k3a [16]),
        .I1(\a7/k4a [16]),
        .O(k6b[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[16]_i_1__6 
       (.I0(\a8/k3a [16]),
        .I1(\a8/k4a [16]),
        .O(k7b[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[16]_i_1__7 
       (.I0(\a9/k3a [16]),
        .I1(\a9/k4a [16]),
        .O(k8b[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[17]_i_1 
       (.I0(\a1/k3a [17]),
        .I1(\a1/k4a [17]),
        .O(k0b[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[17]_i_1__0 
       (.I0(\a2/k3a [17]),
        .I1(\a2/k4a [17]),
        .O(k1b[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[17]_i_1__1 
       (.I0(\a3/k3a [17]),
        .I1(\a3/k4a [17]),
        .O(k2b[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[17]_i_1__2 
       (.I0(\a4/k3a [17]),
        .I1(\a4/k4a [17]),
        .O(k3b[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[17]_i_1__3 
       (.I0(\a5/k3a [17]),
        .I1(\a5/k4a [17]),
        .O(k4b[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[17]_i_1__4 
       (.I0(\a6/k3a [17]),
        .I1(\a6/k4a [17]),
        .O(k5b[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[17]_i_1__5 
       (.I0(\a7/k3a [17]),
        .I1(\a7/k4a [17]),
        .O(k6b[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[17]_i_1__6 
       (.I0(\a8/k3a [17]),
        .I1(\a8/k4a [17]),
        .O(k7b[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[17]_i_1__7 
       (.I0(\a9/k3a [17]),
        .I1(\a9/k4a [17]),
        .O(k8b[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[18]_i_1 
       (.I0(\a1/k3a [18]),
        .I1(\a1/k4a [18]),
        .O(k0b[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[18]_i_1__0 
       (.I0(\a2/k3a [18]),
        .I1(\a2/k4a [18]),
        .O(k1b[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[18]_i_1__1 
       (.I0(\a3/k3a [18]),
        .I1(\a3/k4a [18]),
        .O(k2b[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[18]_i_1__2 
       (.I0(\a4/k3a [18]),
        .I1(\a4/k4a [18]),
        .O(k3b[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[18]_i_1__3 
       (.I0(\a5/k3a [18]),
        .I1(\a5/k4a [18]),
        .O(k4b[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[18]_i_1__4 
       (.I0(\a6/k3a [18]),
        .I1(\a6/k4a [18]),
        .O(k5b[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[18]_i_1__5 
       (.I0(\a7/k3a [18]),
        .I1(\a7/k4a [18]),
        .O(k6b[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[18]_i_1__6 
       (.I0(\a8/k3a [18]),
        .I1(\a8/k4a [18]),
        .O(k7b[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[18]_i_1__7 
       (.I0(\a9/k3a [18]),
        .I1(\a9/k4a [18]),
        .O(k8b[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[19]_i_1 
       (.I0(\a1/k3a [19]),
        .I1(\a1/k4a [19]),
        .O(k0b[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[19]_i_1__0 
       (.I0(\a2/k3a [19]),
        .I1(\a2/k4a [19]),
        .O(k1b[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[19]_i_1__1 
       (.I0(\a3/k3a [19]),
        .I1(\a3/k4a [19]),
        .O(k2b[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[19]_i_1__2 
       (.I0(\a4/k3a [19]),
        .I1(\a4/k4a [19]),
        .O(k3b[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[19]_i_1__3 
       (.I0(\a5/k3a [19]),
        .I1(\a5/k4a [19]),
        .O(k4b[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[19]_i_1__4 
       (.I0(\a6/k3a [19]),
        .I1(\a6/k4a [19]),
        .O(k5b[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[19]_i_1__5 
       (.I0(\a7/k3a [19]),
        .I1(\a7/k4a [19]),
        .O(k6b[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[19]_i_1__6 
       (.I0(\a8/k3a [19]),
        .I1(\a8/k4a [19]),
        .O(k7b[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[19]_i_1__7 
       (.I0(\a9/k3a [19]),
        .I1(\a9/k4a [19]),
        .O(k8b[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[1]_i_1 
       (.I0(\a1/k3a [1]),
        .I1(\a1/k4a [1]),
        .O(k0b[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[1]_i_1__0 
       (.I0(\a2/k3a [1]),
        .I1(\a2/k4a [1]),
        .O(k1b[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[1]_i_1__1 
       (.I0(\a3/k3a [1]),
        .I1(\a3/k4a [1]),
        .O(k2b[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[1]_i_1__2 
       (.I0(\a4/k3a [1]),
        .I1(\a4/k4a [1]),
        .O(k3b[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[1]_i_1__3 
       (.I0(\a5/k3a [1]),
        .I1(\a5/k4a [1]),
        .O(k4b[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[1]_i_1__4 
       (.I0(\a6/k3a [1]),
        .I1(\a6/k4a [1]),
        .O(k5b[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[1]_i_1__5 
       (.I0(\a7/k3a [1]),
        .I1(\a7/k4a [1]),
        .O(k6b[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[1]_i_1__6 
       (.I0(\a8/k3a [1]),
        .I1(\a8/k4a [1]),
        .O(k7b[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[1]_i_1__7 
       (.I0(\a9/k3a [1]),
        .I1(\a9/k4a [1]),
        .O(k8b[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[20]_i_1 
       (.I0(\a1/k3a [20]),
        .I1(\a1/k4a [20]),
        .O(k0b[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[20]_i_1__0 
       (.I0(\a2/k3a [20]),
        .I1(\a2/k4a [20]),
        .O(k1b[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[20]_i_1__1 
       (.I0(\a3/k3a [20]),
        .I1(\a3/k4a [20]),
        .O(k2b[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[20]_i_1__2 
       (.I0(\a4/k3a [20]),
        .I1(\a4/k4a [20]),
        .O(k3b[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[20]_i_1__3 
       (.I0(\a5/k3a [20]),
        .I1(\a5/k4a [20]),
        .O(k4b[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[20]_i_1__4 
       (.I0(\a6/k3a [20]),
        .I1(\a6/k4a [20]),
        .O(k5b[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[20]_i_1__5 
       (.I0(\a7/k3a [20]),
        .I1(\a7/k4a [20]),
        .O(k6b[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[20]_i_1__6 
       (.I0(\a8/k3a [20]),
        .I1(\a8/k4a [20]),
        .O(k7b[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[20]_i_1__7 
       (.I0(\a9/k3a [20]),
        .I1(\a9/k4a [20]),
        .O(k8b[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[21]_i_1 
       (.I0(\a1/k3a [21]),
        .I1(\a1/k4a [21]),
        .O(k0b[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[21]_i_1__0 
       (.I0(\a2/k3a [21]),
        .I1(\a2/k4a [21]),
        .O(k1b[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[21]_i_1__1 
       (.I0(\a3/k3a [21]),
        .I1(\a3/k4a [21]),
        .O(k2b[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[21]_i_1__2 
       (.I0(\a4/k3a [21]),
        .I1(\a4/k4a [21]),
        .O(k3b[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[21]_i_1__3 
       (.I0(\a5/k3a [21]),
        .I1(\a5/k4a [21]),
        .O(k4b[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[21]_i_1__4 
       (.I0(\a6/k3a [21]),
        .I1(\a6/k4a [21]),
        .O(k5b[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[21]_i_1__5 
       (.I0(\a7/k3a [21]),
        .I1(\a7/k4a [21]),
        .O(k6b[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[21]_i_1__6 
       (.I0(\a8/k3a [21]),
        .I1(\a8/k4a [21]),
        .O(k7b[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[21]_i_1__7 
       (.I0(\a9/k3a [21]),
        .I1(\a9/k4a [21]),
        .O(k8b[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[22]_i_1 
       (.I0(\a1/k3a [22]),
        .I1(\a1/k4a [22]),
        .O(k0b[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[22]_i_1__0 
       (.I0(\a2/k3a [22]),
        .I1(\a2/k4a [22]),
        .O(k1b[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[22]_i_1__1 
       (.I0(\a3/k3a [22]),
        .I1(\a3/k4a [22]),
        .O(k2b[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[22]_i_1__2 
       (.I0(\a4/k3a [22]),
        .I1(\a4/k4a [22]),
        .O(k3b[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[22]_i_1__3 
       (.I0(\a5/k3a [22]),
        .I1(\a5/k4a [22]),
        .O(k4b[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[22]_i_1__4 
       (.I0(\a6/k3a [22]),
        .I1(\a6/k4a [22]),
        .O(k5b[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[22]_i_1__5 
       (.I0(\a7/k3a [22]),
        .I1(\a7/k4a [22]),
        .O(k6b[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[22]_i_1__6 
       (.I0(\a8/k3a [22]),
        .I1(\a8/k4a [22]),
        .O(k7b[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[22]_i_1__7 
       (.I0(\a9/k3a [22]),
        .I1(\a9/k4a [22]),
        .O(k8b[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[23]_i_1 
       (.I0(\a1/k3a [23]),
        .I1(\a1/k4a [23]),
        .O(k0b[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[23]_i_1__0 
       (.I0(\a2/k3a [23]),
        .I1(\a2/k4a [23]),
        .O(k1b[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[23]_i_1__1 
       (.I0(\a3/k3a [23]),
        .I1(\a3/k4a [23]),
        .O(k2b[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[23]_i_1__2 
       (.I0(\a4/k3a [23]),
        .I1(\a4/k4a [23]),
        .O(k3b[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[23]_i_1__3 
       (.I0(\a5/k3a [23]),
        .I1(\a5/k4a [23]),
        .O(k4b[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[23]_i_1__4 
       (.I0(\a6/k3a [23]),
        .I1(\a6/k4a [23]),
        .O(k5b[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[23]_i_1__5 
       (.I0(\a7/k3a [23]),
        .I1(\a7/k4a [23]),
        .O(k6b[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[23]_i_1__6 
       (.I0(\a8/k3a [23]),
        .I1(\a8/k4a [23]),
        .O(k7b[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[23]_i_1__7 
       (.I0(\a9/k3a [23]),
        .I1(\a9/k4a [23]),
        .O(k8b[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[24]_i_1 
       (.I0(\a1/k3a [24]),
        .I1(\a1/k4a [24]),
        .O(k0b[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[24]_i_1__0 
       (.I0(\a2/k3a [24]),
        .I1(\a2/k4a [24]),
        .O(k1b[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[24]_i_1__1 
       (.I0(\a3/k3a [24]),
        .I1(\a3/k4a [24]),
        .O(k2b[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[24]_i_1__2 
       (.I0(\a4/k3a [24]),
        .I1(\a4/k4a [24]),
        .O(k3b[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[24]_i_1__3 
       (.I0(\a5/k3a [24]),
        .I1(\a5/k4a [24]),
        .O(k4b[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[24]_i_1__4 
       (.I0(\a6/k3a [24]),
        .I1(\a6/k4a [24]),
        .O(k5b[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[24]_i_1__5 
       (.I0(\a7/k3a [24]),
        .I1(\a7/k4a [24]),
        .O(k6b[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[24]_i_1__6 
       (.I0(\a8/k3a [24]),
        .I1(\a8/k4a [24]),
        .O(k7b[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[24]_i_1__7 
       (.I0(\a9/k3a [24]),
        .I1(\a9/k4a [24]),
        .O(k8b[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[25]_i_1 
       (.I0(\a1/k3a [25]),
        .I1(\a1/k4a [25]),
        .O(k0b[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[25]_i_1__0 
       (.I0(\a2/k3a [25]),
        .I1(\a2/k4a [25]),
        .O(k1b[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[25]_i_1__1 
       (.I0(\a3/k3a [25]),
        .I1(\a3/k4a [25]),
        .O(k2b[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[25]_i_1__2 
       (.I0(\a4/k3a [25]),
        .I1(\a4/k4a [25]),
        .O(k3b[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[25]_i_1__3 
       (.I0(\a5/k3a [25]),
        .I1(\a5/k4a [25]),
        .O(k4b[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[25]_i_1__4 
       (.I0(\a6/k3a [25]),
        .I1(\a6/k4a [25]),
        .O(k5b[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[25]_i_1__5 
       (.I0(\a7/k3a [25]),
        .I1(\a7/k4a [25]),
        .O(k6b[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[25]_i_1__6 
       (.I0(\a8/k3a [25]),
        .I1(\a8/k4a [25]),
        .O(k7b[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[25]_i_1__7 
       (.I0(\a9/k3a [25]),
        .I1(\a9/k4a [25]),
        .O(k8b[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[26]_i_1 
       (.I0(\a1/k3a [26]),
        .I1(\a1/k4a [26]),
        .O(k0b[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[26]_i_1__0 
       (.I0(\a2/k3a [26]),
        .I1(\a2/k4a [26]),
        .O(k1b[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[26]_i_1__1 
       (.I0(\a3/k3a [26]),
        .I1(\a3/k4a [26]),
        .O(k2b[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[26]_i_1__2 
       (.I0(\a4/k3a [26]),
        .I1(\a4/k4a [26]),
        .O(k3b[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[26]_i_1__3 
       (.I0(\a5/k3a [26]),
        .I1(\a5/k4a [26]),
        .O(k4b[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[26]_i_1__4 
       (.I0(\a6/k3a [26]),
        .I1(\a6/k4a [26]),
        .O(k5b[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[26]_i_1__5 
       (.I0(\a7/k3a [26]),
        .I1(\a7/k4a [26]),
        .O(k6b[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[26]_i_1__6 
       (.I0(\a8/k3a [26]),
        .I1(\a8/k4a [26]),
        .O(k7b[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[26]_i_1__7 
       (.I0(\a9/k3a [26]),
        .I1(\a9/k4a [26]),
        .O(k8b[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[27]_i_1 
       (.I0(\a1/k3a [27]),
        .I1(\a1/k4a [27]),
        .O(k0b[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[27]_i_1__0 
       (.I0(\a2/k3a [27]),
        .I1(\a2/k4a [27]),
        .O(k1b[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[27]_i_1__1 
       (.I0(\a3/k3a [27]),
        .I1(\a3/k4a [27]),
        .O(k2b[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[27]_i_1__2 
       (.I0(\a4/k3a [27]),
        .I1(\a4/k4a [27]),
        .O(k3b[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[27]_i_1__3 
       (.I0(\a5/k3a [27]),
        .I1(\a5/k4a [27]),
        .O(k4b[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[27]_i_1__4 
       (.I0(\a6/k3a [27]),
        .I1(\a6/k4a [27]),
        .O(k5b[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[27]_i_1__5 
       (.I0(\a7/k3a [27]),
        .I1(\a7/k4a [27]),
        .O(k6b[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[27]_i_1__6 
       (.I0(\a8/k3a [27]),
        .I1(\a8/k4a [27]),
        .O(k7b[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[27]_i_1__7 
       (.I0(\a9/k3a [27]),
        .I1(\a9/k4a [27]),
        .O(k8b[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[28]_i_1 
       (.I0(\a1/k3a [28]),
        .I1(\a1/k4a [28]),
        .O(k0b[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[28]_i_1__0 
       (.I0(\a2/k3a [28]),
        .I1(\a2/k4a [28]),
        .O(k1b[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[28]_i_1__1 
       (.I0(\a3/k3a [28]),
        .I1(\a3/k4a [28]),
        .O(k2b[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[28]_i_1__2 
       (.I0(\a4/k3a [28]),
        .I1(\a4/k4a [28]),
        .O(k3b[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[28]_i_1__3 
       (.I0(\a5/k3a [28]),
        .I1(\a5/k4a [28]),
        .O(k4b[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[28]_i_1__4 
       (.I0(\a6/k3a [28]),
        .I1(\a6/k4a [28]),
        .O(k5b[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[28]_i_1__5 
       (.I0(\a7/k3a [28]),
        .I1(\a7/k4a [28]),
        .O(k6b[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[28]_i_1__6 
       (.I0(\a8/k3a [28]),
        .I1(\a8/k4a [28]),
        .O(k7b[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[28]_i_1__7 
       (.I0(\a9/k3a [28]),
        .I1(\a9/k4a [28]),
        .O(k8b[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[29]_i_1 
       (.I0(\a1/k3a [29]),
        .I1(\a1/k4a [29]),
        .O(k0b[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[29]_i_1__0 
       (.I0(\a2/k3a [29]),
        .I1(\a2/k4a [29]),
        .O(k1b[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[29]_i_1__1 
       (.I0(\a3/k3a [29]),
        .I1(\a3/k4a [29]),
        .O(k2b[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[29]_i_1__2 
       (.I0(\a4/k3a [29]),
        .I1(\a4/k4a [29]),
        .O(k3b[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[29]_i_1__3 
       (.I0(\a5/k3a [29]),
        .I1(\a5/k4a [29]),
        .O(k4b[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[29]_i_1__4 
       (.I0(\a6/k3a [29]),
        .I1(\a6/k4a [29]),
        .O(k5b[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[29]_i_1__5 
       (.I0(\a7/k3a [29]),
        .I1(\a7/k4a [29]),
        .O(k6b[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[29]_i_1__6 
       (.I0(\a8/k3a [29]),
        .I1(\a8/k4a [29]),
        .O(k7b[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[29]_i_1__7 
       (.I0(\a9/k3a [29]),
        .I1(\a9/k4a [29]),
        .O(k8b[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[2]_i_1 
       (.I0(\a1/k3a [2]),
        .I1(\a1/k4a [2]),
        .O(k0b[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[2]_i_1__0 
       (.I0(\a2/k3a [2]),
        .I1(\a2/k4a [2]),
        .O(k1b[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[2]_i_1__1 
       (.I0(\a3/k3a [2]),
        .I1(\a3/k4a [2]),
        .O(k2b[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[2]_i_1__2 
       (.I0(\a4/k3a [2]),
        .I1(\a4/k4a [2]),
        .O(k3b[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[2]_i_1__3 
       (.I0(\a5/k3a [2]),
        .I1(\a5/k4a [2]),
        .O(k4b[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[2]_i_1__4 
       (.I0(\a6/k3a [2]),
        .I1(\a6/k4a [2]),
        .O(k5b[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[2]_i_1__5 
       (.I0(\a7/k3a [2]),
        .I1(\a7/k4a [2]),
        .O(k6b[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[2]_i_1__6 
       (.I0(\a8/k3a [2]),
        .I1(\a8/k4a [2]),
        .O(k7b[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[2]_i_1__7 
       (.I0(\a9/k3a [2]),
        .I1(\a9/k4a [2]),
        .O(k8b[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[30]_i_1 
       (.I0(\a1/k3a [30]),
        .I1(\a1/k4a [30]),
        .O(k0b[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[30]_i_1__0 
       (.I0(\a2/k3a [30]),
        .I1(\a2/k4a [30]),
        .O(k1b[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[30]_i_1__1 
       (.I0(\a3/k3a [30]),
        .I1(\a3/k4a [30]),
        .O(k2b[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[30]_i_1__2 
       (.I0(\a4/k3a [30]),
        .I1(\a4/k4a [30]),
        .O(k3b[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[30]_i_1__3 
       (.I0(\a5/k3a [30]),
        .I1(\a5/k4a [30]),
        .O(k4b[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[30]_i_1__4 
       (.I0(\a6/k3a [30]),
        .I1(\a6/k4a [30]),
        .O(k5b[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[30]_i_1__5 
       (.I0(\a7/k3a [30]),
        .I1(\a7/k4a [30]),
        .O(k6b[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[30]_i_1__6 
       (.I0(\a8/k3a [30]),
        .I1(\a8/k4a [30]),
        .O(k7b[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[30]_i_1__7 
       (.I0(\a9/k3a [30]),
        .I1(\a9/k4a [30]),
        .O(k8b[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[31]_i_1 
       (.I0(\a1/k3a [31]),
        .I1(\a1/k4a [31]),
        .O(k0b[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[31]_i_1__0 
       (.I0(\a2/k3a [31]),
        .I1(\a2/k4a [31]),
        .O(k1b[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[31]_i_1__1 
       (.I0(\a3/k3a [31]),
        .I1(\a3/k4a [31]),
        .O(k2b[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[31]_i_1__2 
       (.I0(\a4/k3a [31]),
        .I1(\a4/k4a [31]),
        .O(k3b[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[31]_i_1__3 
       (.I0(\a5/k3a [31]),
        .I1(\a5/k4a [31]),
        .O(k4b[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[31]_i_1__4 
       (.I0(\a6/k3a [31]),
        .I1(\a6/k4a [31]),
        .O(k5b[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[31]_i_1__5 
       (.I0(\a7/k3a [31]),
        .I1(\a7/k4a [31]),
        .O(k6b[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[31]_i_1__6 
       (.I0(\a8/k3a [31]),
        .I1(\a8/k4a [31]),
        .O(k7b[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[31]_i_1__7 
       (.I0(\a9/k3a [31]),
        .I1(\a9/k4a [31]),
        .O(k8b[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[32]_i_1 
       (.I0(\a1/k2a [0]),
        .I1(\a1/k4a [0]),
        .O(k0b[32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[32]_i_1__0 
       (.I0(\a2/k2a [0]),
        .I1(\a2/k4a [0]),
        .O(k1b[32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[32]_i_1__1 
       (.I0(\a3/k2a [0]),
        .I1(\a3/k4a [0]),
        .O(k2b[32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[32]_i_1__2 
       (.I0(\a4/k2a [0]),
        .I1(\a4/k4a [0]),
        .O(k3b[32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[32]_i_1__3 
       (.I0(\a5/k2a [0]),
        .I1(\a5/k4a [0]),
        .O(k4b[32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[32]_i_1__4 
       (.I0(\a6/k2a [0]),
        .I1(\a6/k4a [0]),
        .O(k5b[32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[32]_i_1__5 
       (.I0(\a7/k2a [0]),
        .I1(\a7/k4a [0]),
        .O(k6b[32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[32]_i_1__6 
       (.I0(\a8/k2a [0]),
        .I1(\a8/k4a [0]),
        .O(k7b[32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[32]_i_1__7 
       (.I0(\a9/k2a [0]),
        .I1(\a9/k4a [0]),
        .O(k8b[32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[33]_i_1 
       (.I0(\a1/k2a [1]),
        .I1(\a1/k4a [1]),
        .O(k0b[33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[33]_i_1__0 
       (.I0(\a2/k2a [1]),
        .I1(\a2/k4a [1]),
        .O(k1b[33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[33]_i_1__1 
       (.I0(\a3/k2a [1]),
        .I1(\a3/k4a [1]),
        .O(k2b[33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[33]_i_1__2 
       (.I0(\a4/k2a [1]),
        .I1(\a4/k4a [1]),
        .O(k3b[33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[33]_i_1__3 
       (.I0(\a5/k2a [1]),
        .I1(\a5/k4a [1]),
        .O(k4b[33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[33]_i_1__4 
       (.I0(\a6/k2a [1]),
        .I1(\a6/k4a [1]),
        .O(k5b[33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[33]_i_1__5 
       (.I0(\a7/k2a [1]),
        .I1(\a7/k4a [1]),
        .O(k6b[33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[33]_i_1__6 
       (.I0(\a8/k2a [1]),
        .I1(\a8/k4a [1]),
        .O(k7b[33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[33]_i_1__7 
       (.I0(\a9/k2a [1]),
        .I1(\a9/k4a [1]),
        .O(k8b[33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[34]_i_1 
       (.I0(\a1/k2a [2]),
        .I1(\a1/k4a [2]),
        .O(k0b[34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[34]_i_1__0 
       (.I0(\a2/k2a [2]),
        .I1(\a2/k4a [2]),
        .O(k1b[34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[34]_i_1__1 
       (.I0(\a3/k2a [2]),
        .I1(\a3/k4a [2]),
        .O(k2b[34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[34]_i_1__2 
       (.I0(\a4/k2a [2]),
        .I1(\a4/k4a [2]),
        .O(k3b[34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[34]_i_1__3 
       (.I0(\a5/k2a [2]),
        .I1(\a5/k4a [2]),
        .O(k4b[34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[34]_i_1__4 
       (.I0(\a6/k2a [2]),
        .I1(\a6/k4a [2]),
        .O(k5b[34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[34]_i_1__5 
       (.I0(\a7/k2a [2]),
        .I1(\a7/k4a [2]),
        .O(k6b[34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[34]_i_1__6 
       (.I0(\a8/k2a [2]),
        .I1(\a8/k4a [2]),
        .O(k7b[34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[34]_i_1__7 
       (.I0(\a9/k2a [2]),
        .I1(\a9/k4a [2]),
        .O(k8b[34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[35]_i_1 
       (.I0(\a1/k2a [3]),
        .I1(\a1/k4a [3]),
        .O(k0b[35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[35]_i_1__0 
       (.I0(\a2/k2a [3]),
        .I1(\a2/k4a [3]),
        .O(k1b[35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[35]_i_1__1 
       (.I0(\a3/k2a [3]),
        .I1(\a3/k4a [3]),
        .O(k2b[35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[35]_i_1__2 
       (.I0(\a4/k2a [3]),
        .I1(\a4/k4a [3]),
        .O(k3b[35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[35]_i_1__3 
       (.I0(\a5/k2a [3]),
        .I1(\a5/k4a [3]),
        .O(k4b[35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[35]_i_1__4 
       (.I0(\a6/k2a [3]),
        .I1(\a6/k4a [3]),
        .O(k5b[35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[35]_i_1__5 
       (.I0(\a7/k2a [3]),
        .I1(\a7/k4a [3]),
        .O(k6b[35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[35]_i_1__6 
       (.I0(\a8/k2a [3]),
        .I1(\a8/k4a [3]),
        .O(k7b[35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[35]_i_1__7 
       (.I0(\a9/k2a [3]),
        .I1(\a9/k4a [3]),
        .O(k8b[35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[36]_i_1 
       (.I0(\a1/k2a [4]),
        .I1(\a1/k4a [4]),
        .O(k0b[36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[36]_i_1__0 
       (.I0(\a2/k2a [4]),
        .I1(\a2/k4a [4]),
        .O(k1b[36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[36]_i_1__1 
       (.I0(\a3/k2a [4]),
        .I1(\a3/k4a [4]),
        .O(k2b[36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[36]_i_1__2 
       (.I0(\a4/k2a [4]),
        .I1(\a4/k4a [4]),
        .O(k3b[36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[36]_i_1__3 
       (.I0(\a5/k2a [4]),
        .I1(\a5/k4a [4]),
        .O(k4b[36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[36]_i_1__4 
       (.I0(\a6/k2a [4]),
        .I1(\a6/k4a [4]),
        .O(k5b[36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[36]_i_1__5 
       (.I0(\a7/k2a [4]),
        .I1(\a7/k4a [4]),
        .O(k6b[36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[36]_i_1__6 
       (.I0(\a8/k2a [4]),
        .I1(\a8/k4a [4]),
        .O(k7b[36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[36]_i_1__7 
       (.I0(\a9/k2a [4]),
        .I1(\a9/k4a [4]),
        .O(k8b[36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[37]_i_1 
       (.I0(\a1/k2a [5]),
        .I1(\a1/k4a [5]),
        .O(k0b[37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[37]_i_1__0 
       (.I0(\a2/k2a [5]),
        .I1(\a2/k4a [5]),
        .O(k1b[37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[37]_i_1__1 
       (.I0(\a3/k2a [5]),
        .I1(\a3/k4a [5]),
        .O(k2b[37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[37]_i_1__2 
       (.I0(\a4/k2a [5]),
        .I1(\a4/k4a [5]),
        .O(k3b[37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[37]_i_1__3 
       (.I0(\a5/k2a [5]),
        .I1(\a5/k4a [5]),
        .O(k4b[37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[37]_i_1__4 
       (.I0(\a6/k2a [5]),
        .I1(\a6/k4a [5]),
        .O(k5b[37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[37]_i_1__5 
       (.I0(\a7/k2a [5]),
        .I1(\a7/k4a [5]),
        .O(k6b[37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[37]_i_1__6 
       (.I0(\a8/k2a [5]),
        .I1(\a8/k4a [5]),
        .O(k7b[37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[37]_i_1__7 
       (.I0(\a9/k2a [5]),
        .I1(\a9/k4a [5]),
        .O(k8b[37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[38]_i_1 
       (.I0(\a1/k2a [6]),
        .I1(\a1/k4a [6]),
        .O(k0b[38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[38]_i_1__0 
       (.I0(\a2/k2a [6]),
        .I1(\a2/k4a [6]),
        .O(k1b[38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[38]_i_1__1 
       (.I0(\a3/k2a [6]),
        .I1(\a3/k4a [6]),
        .O(k2b[38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[38]_i_1__2 
       (.I0(\a4/k2a [6]),
        .I1(\a4/k4a [6]),
        .O(k3b[38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[38]_i_1__3 
       (.I0(\a5/k2a [6]),
        .I1(\a5/k4a [6]),
        .O(k4b[38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[38]_i_1__4 
       (.I0(\a6/k2a [6]),
        .I1(\a6/k4a [6]),
        .O(k5b[38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[38]_i_1__5 
       (.I0(\a7/k2a [6]),
        .I1(\a7/k4a [6]),
        .O(k6b[38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[38]_i_1__6 
       (.I0(\a8/k2a [6]),
        .I1(\a8/k4a [6]),
        .O(k7b[38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[38]_i_1__7 
       (.I0(\a9/k2a [6]),
        .I1(\a9/k4a [6]),
        .O(k8b[38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[39]_i_1 
       (.I0(\a1/k2a [7]),
        .I1(\a1/k4a [7]),
        .O(k0b[39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[39]_i_1__0 
       (.I0(\a2/k2a [7]),
        .I1(\a2/k4a [7]),
        .O(k1b[39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[39]_i_1__1 
       (.I0(\a3/k2a [7]),
        .I1(\a3/k4a [7]),
        .O(k2b[39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[39]_i_1__2 
       (.I0(\a4/k2a [7]),
        .I1(\a4/k4a [7]),
        .O(k3b[39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[39]_i_1__3 
       (.I0(\a5/k2a [7]),
        .I1(\a5/k4a [7]),
        .O(k4b[39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[39]_i_1__4 
       (.I0(\a6/k2a [7]),
        .I1(\a6/k4a [7]),
        .O(k5b[39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[39]_i_1__5 
       (.I0(\a7/k2a [7]),
        .I1(\a7/k4a [7]),
        .O(k6b[39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[39]_i_1__6 
       (.I0(\a8/k2a [7]),
        .I1(\a8/k4a [7]),
        .O(k7b[39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[39]_i_1__7 
       (.I0(\a9/k2a [7]),
        .I1(\a9/k4a [7]),
        .O(k8b[39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[3]_i_1 
       (.I0(\a1/k3a [3]),
        .I1(\a1/k4a [3]),
        .O(k0b[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[3]_i_1__0 
       (.I0(\a2/k3a [3]),
        .I1(\a2/k4a [3]),
        .O(k1b[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[3]_i_1__1 
       (.I0(\a3/k3a [3]),
        .I1(\a3/k4a [3]),
        .O(k2b[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[3]_i_1__2 
       (.I0(\a4/k3a [3]),
        .I1(\a4/k4a [3]),
        .O(k3b[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[3]_i_1__3 
       (.I0(\a5/k3a [3]),
        .I1(\a5/k4a [3]),
        .O(k4b[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[3]_i_1__4 
       (.I0(\a6/k3a [3]),
        .I1(\a6/k4a [3]),
        .O(k5b[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[3]_i_1__5 
       (.I0(\a7/k3a [3]),
        .I1(\a7/k4a [3]),
        .O(k6b[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[3]_i_1__6 
       (.I0(\a8/k3a [3]),
        .I1(\a8/k4a [3]),
        .O(k7b[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[3]_i_1__7 
       (.I0(\a9/k3a [3]),
        .I1(\a9/k4a [3]),
        .O(k8b[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[40]_i_1 
       (.I0(\a1/k2a [8]),
        .I1(\a1/k4a [8]),
        .O(k0b[40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[40]_i_1__0 
       (.I0(\a2/k2a [8]),
        .I1(\a2/k4a [8]),
        .O(k1b[40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[40]_i_1__1 
       (.I0(\a3/k2a [8]),
        .I1(\a3/k4a [8]),
        .O(k2b[40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[40]_i_1__2 
       (.I0(\a4/k2a [8]),
        .I1(\a4/k4a [8]),
        .O(k3b[40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[40]_i_1__3 
       (.I0(\a5/k2a [8]),
        .I1(\a5/k4a [8]),
        .O(k4b[40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[40]_i_1__4 
       (.I0(\a6/k2a [8]),
        .I1(\a6/k4a [8]),
        .O(k5b[40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[40]_i_1__5 
       (.I0(\a7/k2a [8]),
        .I1(\a7/k4a [8]),
        .O(k6b[40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[40]_i_1__6 
       (.I0(\a8/k2a [8]),
        .I1(\a8/k4a [8]),
        .O(k7b[40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[40]_i_1__7 
       (.I0(\a9/k2a [8]),
        .I1(\a9/k4a [8]),
        .O(k8b[40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[41]_i_1 
       (.I0(\a1/k2a [9]),
        .I1(\a1/k4a [9]),
        .O(k0b[41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[41]_i_1__0 
       (.I0(\a2/k2a [9]),
        .I1(\a2/k4a [9]),
        .O(k1b[41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[41]_i_1__1 
       (.I0(\a3/k2a [9]),
        .I1(\a3/k4a [9]),
        .O(k2b[41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[41]_i_1__2 
       (.I0(\a4/k2a [9]),
        .I1(\a4/k4a [9]),
        .O(k3b[41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[41]_i_1__3 
       (.I0(\a5/k2a [9]),
        .I1(\a5/k4a [9]),
        .O(k4b[41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[41]_i_1__4 
       (.I0(\a6/k2a [9]),
        .I1(\a6/k4a [9]),
        .O(k5b[41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[41]_i_1__5 
       (.I0(\a7/k2a [9]),
        .I1(\a7/k4a [9]),
        .O(k6b[41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[41]_i_1__6 
       (.I0(\a8/k2a [9]),
        .I1(\a8/k4a [9]),
        .O(k7b[41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[41]_i_1__7 
       (.I0(\a9/k2a [9]),
        .I1(\a9/k4a [9]),
        .O(k8b[41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[42]_i_1 
       (.I0(\a1/k2a [10]),
        .I1(\a1/k4a [10]),
        .O(k0b[42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[42]_i_1__0 
       (.I0(\a2/k2a [10]),
        .I1(\a2/k4a [10]),
        .O(k1b[42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[42]_i_1__1 
       (.I0(\a3/k2a [10]),
        .I1(\a3/k4a [10]),
        .O(k2b[42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[42]_i_1__2 
       (.I0(\a4/k2a [10]),
        .I1(\a4/k4a [10]),
        .O(k3b[42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[42]_i_1__3 
       (.I0(\a5/k2a [10]),
        .I1(\a5/k4a [10]),
        .O(k4b[42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[42]_i_1__4 
       (.I0(\a6/k2a [10]),
        .I1(\a6/k4a [10]),
        .O(k5b[42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[42]_i_1__5 
       (.I0(\a7/k2a [10]),
        .I1(\a7/k4a [10]),
        .O(k6b[42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[42]_i_1__6 
       (.I0(\a8/k2a [10]),
        .I1(\a8/k4a [10]),
        .O(k7b[42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[42]_i_1__7 
       (.I0(\a9/k2a [10]),
        .I1(\a9/k4a [10]),
        .O(k8b[42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[43]_i_1 
       (.I0(\a1/k2a [11]),
        .I1(\a1/k4a [11]),
        .O(k0b[43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[43]_i_1__0 
       (.I0(\a2/k2a [11]),
        .I1(\a2/k4a [11]),
        .O(k1b[43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[43]_i_1__1 
       (.I0(\a3/k2a [11]),
        .I1(\a3/k4a [11]),
        .O(k2b[43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[43]_i_1__2 
       (.I0(\a4/k2a [11]),
        .I1(\a4/k4a [11]),
        .O(k3b[43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[43]_i_1__3 
       (.I0(\a5/k2a [11]),
        .I1(\a5/k4a [11]),
        .O(k4b[43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[43]_i_1__4 
       (.I0(\a6/k2a [11]),
        .I1(\a6/k4a [11]),
        .O(k5b[43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[43]_i_1__5 
       (.I0(\a7/k2a [11]),
        .I1(\a7/k4a [11]),
        .O(k6b[43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[43]_i_1__6 
       (.I0(\a8/k2a [11]),
        .I1(\a8/k4a [11]),
        .O(k7b[43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[43]_i_1__7 
       (.I0(\a9/k2a [11]),
        .I1(\a9/k4a [11]),
        .O(k8b[43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[44]_i_1 
       (.I0(\a1/k2a [12]),
        .I1(\a1/k4a [12]),
        .O(k0b[44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[44]_i_1__0 
       (.I0(\a2/k2a [12]),
        .I1(\a2/k4a [12]),
        .O(k1b[44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[44]_i_1__1 
       (.I0(\a3/k2a [12]),
        .I1(\a3/k4a [12]),
        .O(k2b[44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[44]_i_1__2 
       (.I0(\a4/k2a [12]),
        .I1(\a4/k4a [12]),
        .O(k3b[44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[44]_i_1__3 
       (.I0(\a5/k2a [12]),
        .I1(\a5/k4a [12]),
        .O(k4b[44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[44]_i_1__4 
       (.I0(\a6/k2a [12]),
        .I1(\a6/k4a [12]),
        .O(k5b[44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[44]_i_1__5 
       (.I0(\a7/k2a [12]),
        .I1(\a7/k4a [12]),
        .O(k6b[44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[44]_i_1__6 
       (.I0(\a8/k2a [12]),
        .I1(\a8/k4a [12]),
        .O(k7b[44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[44]_i_1__7 
       (.I0(\a9/k2a [12]),
        .I1(\a9/k4a [12]),
        .O(k8b[44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[45]_i_1 
       (.I0(\a1/k2a [13]),
        .I1(\a1/k4a [13]),
        .O(k0b[45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[45]_i_1__0 
       (.I0(\a2/k2a [13]),
        .I1(\a2/k4a [13]),
        .O(k1b[45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[45]_i_1__1 
       (.I0(\a3/k2a [13]),
        .I1(\a3/k4a [13]),
        .O(k2b[45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[45]_i_1__2 
       (.I0(\a4/k2a [13]),
        .I1(\a4/k4a [13]),
        .O(k3b[45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[45]_i_1__3 
       (.I0(\a5/k2a [13]),
        .I1(\a5/k4a [13]),
        .O(k4b[45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[45]_i_1__4 
       (.I0(\a6/k2a [13]),
        .I1(\a6/k4a [13]),
        .O(k5b[45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[45]_i_1__5 
       (.I0(\a7/k2a [13]),
        .I1(\a7/k4a [13]),
        .O(k6b[45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[45]_i_1__6 
       (.I0(\a8/k2a [13]),
        .I1(\a8/k4a [13]),
        .O(k7b[45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[45]_i_1__7 
       (.I0(\a9/k2a [13]),
        .I1(\a9/k4a [13]),
        .O(k8b[45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[46]_i_1 
       (.I0(\a1/k2a [14]),
        .I1(\a1/k4a [14]),
        .O(k0b[46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[46]_i_1__0 
       (.I0(\a2/k2a [14]),
        .I1(\a2/k4a [14]),
        .O(k1b[46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[46]_i_1__1 
       (.I0(\a3/k2a [14]),
        .I1(\a3/k4a [14]),
        .O(k2b[46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[46]_i_1__2 
       (.I0(\a4/k2a [14]),
        .I1(\a4/k4a [14]),
        .O(k3b[46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[46]_i_1__3 
       (.I0(\a5/k2a [14]),
        .I1(\a5/k4a [14]),
        .O(k4b[46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[46]_i_1__4 
       (.I0(\a6/k2a [14]),
        .I1(\a6/k4a [14]),
        .O(k5b[46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[46]_i_1__5 
       (.I0(\a7/k2a [14]),
        .I1(\a7/k4a [14]),
        .O(k6b[46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[46]_i_1__6 
       (.I0(\a8/k2a [14]),
        .I1(\a8/k4a [14]),
        .O(k7b[46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[46]_i_1__7 
       (.I0(\a9/k2a [14]),
        .I1(\a9/k4a [14]),
        .O(k8b[46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[47]_i_1 
       (.I0(\a1/k2a [15]),
        .I1(\a1/k4a [15]),
        .O(k0b[47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[47]_i_1__0 
       (.I0(\a2/k2a [15]),
        .I1(\a2/k4a [15]),
        .O(k1b[47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[47]_i_1__1 
       (.I0(\a3/k2a [15]),
        .I1(\a3/k4a [15]),
        .O(k2b[47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[47]_i_1__2 
       (.I0(\a4/k2a [15]),
        .I1(\a4/k4a [15]),
        .O(k3b[47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[47]_i_1__3 
       (.I0(\a5/k2a [15]),
        .I1(\a5/k4a [15]),
        .O(k4b[47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[47]_i_1__4 
       (.I0(\a6/k2a [15]),
        .I1(\a6/k4a [15]),
        .O(k5b[47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[47]_i_1__5 
       (.I0(\a7/k2a [15]),
        .I1(\a7/k4a [15]),
        .O(k6b[47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[47]_i_1__6 
       (.I0(\a8/k2a [15]),
        .I1(\a8/k4a [15]),
        .O(k7b[47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[47]_i_1__7 
       (.I0(\a9/k2a [15]),
        .I1(\a9/k4a [15]),
        .O(k8b[47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[48]_i_1 
       (.I0(\a1/k2a [16]),
        .I1(\a1/k4a [16]),
        .O(k0b[48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[48]_i_1__0 
       (.I0(\a2/k2a [16]),
        .I1(\a2/k4a [16]),
        .O(k1b[48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[48]_i_1__1 
       (.I0(\a3/k2a [16]),
        .I1(\a3/k4a [16]),
        .O(k2b[48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[48]_i_1__2 
       (.I0(\a4/k2a [16]),
        .I1(\a4/k4a [16]),
        .O(k3b[48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[48]_i_1__3 
       (.I0(\a5/k2a [16]),
        .I1(\a5/k4a [16]),
        .O(k4b[48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[48]_i_1__4 
       (.I0(\a6/k2a [16]),
        .I1(\a6/k4a [16]),
        .O(k5b[48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[48]_i_1__5 
       (.I0(\a7/k2a [16]),
        .I1(\a7/k4a [16]),
        .O(k6b[48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[48]_i_1__6 
       (.I0(\a8/k2a [16]),
        .I1(\a8/k4a [16]),
        .O(k7b[48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[48]_i_1__7 
       (.I0(\a9/k2a [16]),
        .I1(\a9/k4a [16]),
        .O(k8b[48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[49]_i_1 
       (.I0(\a1/k2a [17]),
        .I1(\a1/k4a [17]),
        .O(k0b[49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[49]_i_1__0 
       (.I0(\a2/k2a [17]),
        .I1(\a2/k4a [17]),
        .O(k1b[49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[49]_i_1__1 
       (.I0(\a3/k2a [17]),
        .I1(\a3/k4a [17]),
        .O(k2b[49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[49]_i_1__2 
       (.I0(\a4/k2a [17]),
        .I1(\a4/k4a [17]),
        .O(k3b[49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[49]_i_1__3 
       (.I0(\a5/k2a [17]),
        .I1(\a5/k4a [17]),
        .O(k4b[49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[49]_i_1__4 
       (.I0(\a6/k2a [17]),
        .I1(\a6/k4a [17]),
        .O(k5b[49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[49]_i_1__5 
       (.I0(\a7/k2a [17]),
        .I1(\a7/k4a [17]),
        .O(k6b[49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[49]_i_1__6 
       (.I0(\a8/k2a [17]),
        .I1(\a8/k4a [17]),
        .O(k7b[49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[49]_i_1__7 
       (.I0(\a9/k2a [17]),
        .I1(\a9/k4a [17]),
        .O(k8b[49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[4]_i_1 
       (.I0(\a1/k3a [4]),
        .I1(\a1/k4a [4]),
        .O(k0b[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[4]_i_1__0 
       (.I0(\a2/k3a [4]),
        .I1(\a2/k4a [4]),
        .O(k1b[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[4]_i_1__1 
       (.I0(\a3/k3a [4]),
        .I1(\a3/k4a [4]),
        .O(k2b[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[4]_i_1__2 
       (.I0(\a4/k3a [4]),
        .I1(\a4/k4a [4]),
        .O(k3b[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[4]_i_1__3 
       (.I0(\a5/k3a [4]),
        .I1(\a5/k4a [4]),
        .O(k4b[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[4]_i_1__4 
       (.I0(\a6/k3a [4]),
        .I1(\a6/k4a [4]),
        .O(k5b[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[4]_i_1__5 
       (.I0(\a7/k3a [4]),
        .I1(\a7/k4a [4]),
        .O(k6b[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[4]_i_1__6 
       (.I0(\a8/k3a [4]),
        .I1(\a8/k4a [4]),
        .O(k7b[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[4]_i_1__7 
       (.I0(\a9/k3a [4]),
        .I1(\a9/k4a [4]),
        .O(k8b[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[50]_i_1 
       (.I0(\a1/k2a [18]),
        .I1(\a1/k4a [18]),
        .O(k0b[50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[50]_i_1__0 
       (.I0(\a2/k2a [18]),
        .I1(\a2/k4a [18]),
        .O(k1b[50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[50]_i_1__1 
       (.I0(\a3/k2a [18]),
        .I1(\a3/k4a [18]),
        .O(k2b[50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[50]_i_1__2 
       (.I0(\a4/k2a [18]),
        .I1(\a4/k4a [18]),
        .O(k3b[50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[50]_i_1__3 
       (.I0(\a5/k2a [18]),
        .I1(\a5/k4a [18]),
        .O(k4b[50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[50]_i_1__4 
       (.I0(\a6/k2a [18]),
        .I1(\a6/k4a [18]),
        .O(k5b[50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[50]_i_1__5 
       (.I0(\a7/k2a [18]),
        .I1(\a7/k4a [18]),
        .O(k6b[50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[50]_i_1__6 
       (.I0(\a8/k2a [18]),
        .I1(\a8/k4a [18]),
        .O(k7b[50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[50]_i_1__7 
       (.I0(\a9/k2a [18]),
        .I1(\a9/k4a [18]),
        .O(k8b[50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[51]_i_1 
       (.I0(\a1/k2a [19]),
        .I1(\a1/k4a [19]),
        .O(k0b[51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[51]_i_1__0 
       (.I0(\a2/k2a [19]),
        .I1(\a2/k4a [19]),
        .O(k1b[51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[51]_i_1__1 
       (.I0(\a3/k2a [19]),
        .I1(\a3/k4a [19]),
        .O(k2b[51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[51]_i_1__2 
       (.I0(\a4/k2a [19]),
        .I1(\a4/k4a [19]),
        .O(k3b[51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[51]_i_1__3 
       (.I0(\a5/k2a [19]),
        .I1(\a5/k4a [19]),
        .O(k4b[51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[51]_i_1__4 
       (.I0(\a6/k2a [19]),
        .I1(\a6/k4a [19]),
        .O(k5b[51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[51]_i_1__5 
       (.I0(\a7/k2a [19]),
        .I1(\a7/k4a [19]),
        .O(k6b[51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[51]_i_1__6 
       (.I0(\a8/k2a [19]),
        .I1(\a8/k4a [19]),
        .O(k7b[51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[51]_i_1__7 
       (.I0(\a9/k2a [19]),
        .I1(\a9/k4a [19]),
        .O(k8b[51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[52]_i_1 
       (.I0(\a1/k2a [20]),
        .I1(\a1/k4a [20]),
        .O(k0b[52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[52]_i_1__0 
       (.I0(\a2/k2a [20]),
        .I1(\a2/k4a [20]),
        .O(k1b[52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[52]_i_1__1 
       (.I0(\a3/k2a [20]),
        .I1(\a3/k4a [20]),
        .O(k2b[52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[52]_i_1__2 
       (.I0(\a4/k2a [20]),
        .I1(\a4/k4a [20]),
        .O(k3b[52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[52]_i_1__3 
       (.I0(\a5/k2a [20]),
        .I1(\a5/k4a [20]),
        .O(k4b[52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[52]_i_1__4 
       (.I0(\a6/k2a [20]),
        .I1(\a6/k4a [20]),
        .O(k5b[52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[52]_i_1__5 
       (.I0(\a7/k2a [20]),
        .I1(\a7/k4a [20]),
        .O(k6b[52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[52]_i_1__6 
       (.I0(\a8/k2a [20]),
        .I1(\a8/k4a [20]),
        .O(k7b[52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[52]_i_1__7 
       (.I0(\a9/k2a [20]),
        .I1(\a9/k4a [20]),
        .O(k8b[52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[53]_i_1 
       (.I0(\a1/k2a [21]),
        .I1(\a1/k4a [21]),
        .O(k0b[53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[53]_i_1__0 
       (.I0(\a2/k2a [21]),
        .I1(\a2/k4a [21]),
        .O(k1b[53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[53]_i_1__1 
       (.I0(\a3/k2a [21]),
        .I1(\a3/k4a [21]),
        .O(k2b[53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[53]_i_1__2 
       (.I0(\a4/k2a [21]),
        .I1(\a4/k4a [21]),
        .O(k3b[53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[53]_i_1__3 
       (.I0(\a5/k2a [21]),
        .I1(\a5/k4a [21]),
        .O(k4b[53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[53]_i_1__4 
       (.I0(\a6/k2a [21]),
        .I1(\a6/k4a [21]),
        .O(k5b[53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[53]_i_1__5 
       (.I0(\a7/k2a [21]),
        .I1(\a7/k4a [21]),
        .O(k6b[53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[53]_i_1__6 
       (.I0(\a8/k2a [21]),
        .I1(\a8/k4a [21]),
        .O(k7b[53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[53]_i_1__7 
       (.I0(\a9/k2a [21]),
        .I1(\a9/k4a [21]),
        .O(k8b[53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[54]_i_1 
       (.I0(\a1/k2a [22]),
        .I1(\a1/k4a [22]),
        .O(k0b[54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[54]_i_1__0 
       (.I0(\a2/k2a [22]),
        .I1(\a2/k4a [22]),
        .O(k1b[54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[54]_i_1__1 
       (.I0(\a3/k2a [22]),
        .I1(\a3/k4a [22]),
        .O(k2b[54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[54]_i_1__2 
       (.I0(\a4/k2a [22]),
        .I1(\a4/k4a [22]),
        .O(k3b[54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[54]_i_1__3 
       (.I0(\a5/k2a [22]),
        .I1(\a5/k4a [22]),
        .O(k4b[54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[54]_i_1__4 
       (.I0(\a6/k2a [22]),
        .I1(\a6/k4a [22]),
        .O(k5b[54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[54]_i_1__5 
       (.I0(\a7/k2a [22]),
        .I1(\a7/k4a [22]),
        .O(k6b[54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[54]_i_1__6 
       (.I0(\a8/k2a [22]),
        .I1(\a8/k4a [22]),
        .O(k7b[54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[54]_i_1__7 
       (.I0(\a9/k2a [22]),
        .I1(\a9/k4a [22]),
        .O(k8b[54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[55]_i_1 
       (.I0(\a1/k2a [23]),
        .I1(\a1/k4a [23]),
        .O(k0b[55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[55]_i_1__0 
       (.I0(\a2/k2a [23]),
        .I1(\a2/k4a [23]),
        .O(k1b[55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[55]_i_1__1 
       (.I0(\a3/k2a [23]),
        .I1(\a3/k4a [23]),
        .O(k2b[55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[55]_i_1__2 
       (.I0(\a4/k2a [23]),
        .I1(\a4/k4a [23]),
        .O(k3b[55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[55]_i_1__3 
       (.I0(\a5/k2a [23]),
        .I1(\a5/k4a [23]),
        .O(k4b[55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[55]_i_1__4 
       (.I0(\a6/k2a [23]),
        .I1(\a6/k4a [23]),
        .O(k5b[55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[55]_i_1__5 
       (.I0(\a7/k2a [23]),
        .I1(\a7/k4a [23]),
        .O(k6b[55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[55]_i_1__6 
       (.I0(\a8/k2a [23]),
        .I1(\a8/k4a [23]),
        .O(k7b[55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[55]_i_1__7 
       (.I0(\a9/k2a [23]),
        .I1(\a9/k4a [23]),
        .O(k8b[55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[56]_i_1 
       (.I0(\a1/k2a [24]),
        .I1(\a1/k4a [24]),
        .O(k0b[56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[56]_i_1__0 
       (.I0(\a2/k2a [24]),
        .I1(\a2/k4a [24]),
        .O(k1b[56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[56]_i_1__1 
       (.I0(\a3/k2a [24]),
        .I1(\a3/k4a [24]),
        .O(k2b[56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[56]_i_1__2 
       (.I0(\a4/k2a [24]),
        .I1(\a4/k4a [24]),
        .O(k3b[56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[56]_i_1__3 
       (.I0(\a5/k2a [24]),
        .I1(\a5/k4a [24]),
        .O(k4b[56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[56]_i_1__4 
       (.I0(\a6/k2a [24]),
        .I1(\a6/k4a [24]),
        .O(k5b[56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[56]_i_1__5 
       (.I0(\a7/k2a [24]),
        .I1(\a7/k4a [24]),
        .O(k6b[56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[56]_i_1__6 
       (.I0(\a8/k2a [24]),
        .I1(\a8/k4a [24]),
        .O(k7b[56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[56]_i_1__7 
       (.I0(\a9/k2a [24]),
        .I1(\a9/k4a [24]),
        .O(k8b[56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[57]_i_1 
       (.I0(\a1/k2a [25]),
        .I1(\a1/k4a [25]),
        .O(k0b[57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[57]_i_1__0 
       (.I0(\a2/k2a [25]),
        .I1(\a2/k4a [25]),
        .O(k1b[57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[57]_i_1__1 
       (.I0(\a3/k2a [25]),
        .I1(\a3/k4a [25]),
        .O(k2b[57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[57]_i_1__2 
       (.I0(\a4/k2a [25]),
        .I1(\a4/k4a [25]),
        .O(k3b[57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[57]_i_1__3 
       (.I0(\a5/k2a [25]),
        .I1(\a5/k4a [25]),
        .O(k4b[57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[57]_i_1__4 
       (.I0(\a6/k2a [25]),
        .I1(\a6/k4a [25]),
        .O(k5b[57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[57]_i_1__5 
       (.I0(\a7/k2a [25]),
        .I1(\a7/k4a [25]),
        .O(k6b[57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[57]_i_1__6 
       (.I0(\a8/k2a [25]),
        .I1(\a8/k4a [25]),
        .O(k7b[57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[57]_i_1__7 
       (.I0(\a9/k2a [25]),
        .I1(\a9/k4a [25]),
        .O(k8b[57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[58]_i_1 
       (.I0(\a1/k2a [26]),
        .I1(\a1/k4a [26]),
        .O(k0b[58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[58]_i_1__0 
       (.I0(\a2/k2a [26]),
        .I1(\a2/k4a [26]),
        .O(k1b[58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[58]_i_1__1 
       (.I0(\a3/k2a [26]),
        .I1(\a3/k4a [26]),
        .O(k2b[58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[58]_i_1__2 
       (.I0(\a4/k2a [26]),
        .I1(\a4/k4a [26]),
        .O(k3b[58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[58]_i_1__3 
       (.I0(\a5/k2a [26]),
        .I1(\a5/k4a [26]),
        .O(k4b[58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[58]_i_1__4 
       (.I0(\a6/k2a [26]),
        .I1(\a6/k4a [26]),
        .O(k5b[58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[58]_i_1__5 
       (.I0(\a7/k2a [26]),
        .I1(\a7/k4a [26]),
        .O(k6b[58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[58]_i_1__6 
       (.I0(\a8/k2a [26]),
        .I1(\a8/k4a [26]),
        .O(k7b[58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[58]_i_1__7 
       (.I0(\a9/k2a [26]),
        .I1(\a9/k4a [26]),
        .O(k8b[58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[59]_i_1 
       (.I0(\a1/k2a [27]),
        .I1(\a1/k4a [27]),
        .O(k0b[59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[59]_i_1__0 
       (.I0(\a2/k2a [27]),
        .I1(\a2/k4a [27]),
        .O(k1b[59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[59]_i_1__1 
       (.I0(\a3/k2a [27]),
        .I1(\a3/k4a [27]),
        .O(k2b[59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[59]_i_1__2 
       (.I0(\a4/k2a [27]),
        .I1(\a4/k4a [27]),
        .O(k3b[59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[59]_i_1__3 
       (.I0(\a5/k2a [27]),
        .I1(\a5/k4a [27]),
        .O(k4b[59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[59]_i_1__4 
       (.I0(\a6/k2a [27]),
        .I1(\a6/k4a [27]),
        .O(k5b[59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[59]_i_1__5 
       (.I0(\a7/k2a [27]),
        .I1(\a7/k4a [27]),
        .O(k6b[59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[59]_i_1__6 
       (.I0(\a8/k2a [27]),
        .I1(\a8/k4a [27]),
        .O(k7b[59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[59]_i_1__7 
       (.I0(\a9/k2a [27]),
        .I1(\a9/k4a [27]),
        .O(k8b[59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[5]_i_1 
       (.I0(\a1/k3a [5]),
        .I1(\a1/k4a [5]),
        .O(k0b[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[5]_i_1__0 
       (.I0(\a2/k3a [5]),
        .I1(\a2/k4a [5]),
        .O(k1b[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[5]_i_1__1 
       (.I0(\a3/k3a [5]),
        .I1(\a3/k4a [5]),
        .O(k2b[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[5]_i_1__2 
       (.I0(\a4/k3a [5]),
        .I1(\a4/k4a [5]),
        .O(k3b[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[5]_i_1__3 
       (.I0(\a5/k3a [5]),
        .I1(\a5/k4a [5]),
        .O(k4b[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[5]_i_1__4 
       (.I0(\a6/k3a [5]),
        .I1(\a6/k4a [5]),
        .O(k5b[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[5]_i_1__5 
       (.I0(\a7/k3a [5]),
        .I1(\a7/k4a [5]),
        .O(k6b[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[5]_i_1__6 
       (.I0(\a8/k3a [5]),
        .I1(\a8/k4a [5]),
        .O(k7b[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[5]_i_1__7 
       (.I0(\a9/k3a [5]),
        .I1(\a9/k4a [5]),
        .O(k8b[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[60]_i_1 
       (.I0(\a1/k2a [28]),
        .I1(\a1/k4a [28]),
        .O(k0b[60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[60]_i_1__0 
       (.I0(\a2/k2a [28]),
        .I1(\a2/k4a [28]),
        .O(k1b[60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[60]_i_1__1 
       (.I0(\a3/k2a [28]),
        .I1(\a3/k4a [28]),
        .O(k2b[60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[60]_i_1__2 
       (.I0(\a4/k2a [28]),
        .I1(\a4/k4a [28]),
        .O(k3b[60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[60]_i_1__3 
       (.I0(\a5/k2a [28]),
        .I1(\a5/k4a [28]),
        .O(k4b[60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[60]_i_1__4 
       (.I0(\a6/k2a [28]),
        .I1(\a6/k4a [28]),
        .O(k5b[60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[60]_i_1__5 
       (.I0(\a7/k2a [28]),
        .I1(\a7/k4a [28]),
        .O(k6b[60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[60]_i_1__6 
       (.I0(\a8/k2a [28]),
        .I1(\a8/k4a [28]),
        .O(k7b[60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[60]_i_1__7 
       (.I0(\a9/k2a [28]),
        .I1(\a9/k4a [28]),
        .O(k8b[60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[61]_i_1 
       (.I0(\a1/k2a [29]),
        .I1(\a1/k4a [29]),
        .O(k0b[61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[61]_i_1__0 
       (.I0(\a2/k2a [29]),
        .I1(\a2/k4a [29]),
        .O(k1b[61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[61]_i_1__1 
       (.I0(\a3/k2a [29]),
        .I1(\a3/k4a [29]),
        .O(k2b[61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[61]_i_1__2 
       (.I0(\a4/k2a [29]),
        .I1(\a4/k4a [29]),
        .O(k3b[61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[61]_i_1__3 
       (.I0(\a5/k2a [29]),
        .I1(\a5/k4a [29]),
        .O(k4b[61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[61]_i_1__4 
       (.I0(\a6/k2a [29]),
        .I1(\a6/k4a [29]),
        .O(k5b[61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[61]_i_1__5 
       (.I0(\a7/k2a [29]),
        .I1(\a7/k4a [29]),
        .O(k6b[61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[61]_i_1__6 
       (.I0(\a8/k2a [29]),
        .I1(\a8/k4a [29]),
        .O(k7b[61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[61]_i_1__7 
       (.I0(\a9/k2a [29]),
        .I1(\a9/k4a [29]),
        .O(k8b[61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[62]_i_1 
       (.I0(\a1/k2a [30]),
        .I1(\a1/k4a [30]),
        .O(k0b[62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[62]_i_1__0 
       (.I0(\a2/k2a [30]),
        .I1(\a2/k4a [30]),
        .O(k1b[62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[62]_i_1__1 
       (.I0(\a3/k2a [30]),
        .I1(\a3/k4a [30]),
        .O(k2b[62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[62]_i_1__2 
       (.I0(\a4/k2a [30]),
        .I1(\a4/k4a [30]),
        .O(k3b[62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[62]_i_1__3 
       (.I0(\a5/k2a [30]),
        .I1(\a5/k4a [30]),
        .O(k4b[62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[62]_i_1__4 
       (.I0(\a6/k2a [30]),
        .I1(\a6/k4a [30]),
        .O(k5b[62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[62]_i_1__5 
       (.I0(\a7/k2a [30]),
        .I1(\a7/k4a [30]),
        .O(k6b[62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[62]_i_1__6 
       (.I0(\a8/k2a [30]),
        .I1(\a8/k4a [30]),
        .O(k7b[62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[62]_i_1__7 
       (.I0(\a9/k2a [30]),
        .I1(\a9/k4a [30]),
        .O(k8b[62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[63]_i_1 
       (.I0(\a1/k2a [31]),
        .I1(\a1/k4a [31]),
        .O(k0b[63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[63]_i_1__0 
       (.I0(\a2/k2a [31]),
        .I1(\a2/k4a [31]),
        .O(k1b[63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[63]_i_1__1 
       (.I0(\a3/k2a [31]),
        .I1(\a3/k4a [31]),
        .O(k2b[63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[63]_i_1__2 
       (.I0(\a4/k2a [31]),
        .I1(\a4/k4a [31]),
        .O(k3b[63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[63]_i_1__3 
       (.I0(\a5/k2a [31]),
        .I1(\a5/k4a [31]),
        .O(k4b[63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[63]_i_1__4 
       (.I0(\a6/k2a [31]),
        .I1(\a6/k4a [31]),
        .O(k5b[63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[63]_i_1__5 
       (.I0(\a7/k2a [31]),
        .I1(\a7/k4a [31]),
        .O(k6b[63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[63]_i_1__6 
       (.I0(\a8/k2a [31]),
        .I1(\a8/k4a [31]),
        .O(k7b[63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[63]_i_1__7 
       (.I0(\a9/k2a [31]),
        .I1(\a9/k4a [31]),
        .O(k8b[63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[64]_i_1 
       (.I0(\a1/k1a [0]),
        .I1(\a1/k4a [0]),
        .O(k0b[64]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[64]_i_1__0 
       (.I0(\a2/k1a [0]),
        .I1(\a2/k4a [0]),
        .O(k1b[64]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[64]_i_1__1 
       (.I0(\a3/k1a [0]),
        .I1(\a3/k4a [0]),
        .O(k2b[64]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[64]_i_1__2 
       (.I0(\a4/k1a [0]),
        .I1(\a4/k4a [0]),
        .O(k3b[64]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[64]_i_1__3 
       (.I0(\a5/k1a [0]),
        .I1(\a5/k4a [0]),
        .O(k4b[64]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[64]_i_1__4 
       (.I0(\a6/k1a [0]),
        .I1(\a6/k4a [0]),
        .O(k5b[64]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[64]_i_1__5 
       (.I0(\a7/k1a [0]),
        .I1(\a7/k4a [0]),
        .O(k6b[64]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[64]_i_1__6 
       (.I0(\a8/k1a [0]),
        .I1(\a8/k4a [0]),
        .O(k7b[64]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[64]_i_1__7 
       (.I0(\a9/k1a [0]),
        .I1(\a9/k4a [0]),
        .O(k8b[64]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[65]_i_1 
       (.I0(\a1/k1a [1]),
        .I1(\a1/k4a [1]),
        .O(k0b[65]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[65]_i_1__0 
       (.I0(\a2/k1a [1]),
        .I1(\a2/k4a [1]),
        .O(k1b[65]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[65]_i_1__1 
       (.I0(\a3/k1a [1]),
        .I1(\a3/k4a [1]),
        .O(k2b[65]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[65]_i_1__2 
       (.I0(\a4/k1a [1]),
        .I1(\a4/k4a [1]),
        .O(k3b[65]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[65]_i_1__3 
       (.I0(\a5/k1a [1]),
        .I1(\a5/k4a [1]),
        .O(k4b[65]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[65]_i_1__4 
       (.I0(\a6/k1a [1]),
        .I1(\a6/k4a [1]),
        .O(k5b[65]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[65]_i_1__5 
       (.I0(\a7/k1a [1]),
        .I1(\a7/k4a [1]),
        .O(k6b[65]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[65]_i_1__6 
       (.I0(\a8/k1a [1]),
        .I1(\a8/k4a [1]),
        .O(k7b[65]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[65]_i_1__7 
       (.I0(\a9/k1a [1]),
        .I1(\a9/k4a [1]),
        .O(k8b[65]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[66]_i_1 
       (.I0(\a1/k1a [2]),
        .I1(\a1/k4a [2]),
        .O(k0b[66]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[66]_i_1__0 
       (.I0(\a2/k1a [2]),
        .I1(\a2/k4a [2]),
        .O(k1b[66]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[66]_i_1__1 
       (.I0(\a3/k1a [2]),
        .I1(\a3/k4a [2]),
        .O(k2b[66]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[66]_i_1__2 
       (.I0(\a4/k1a [2]),
        .I1(\a4/k4a [2]),
        .O(k3b[66]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[66]_i_1__3 
       (.I0(\a5/k1a [2]),
        .I1(\a5/k4a [2]),
        .O(k4b[66]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[66]_i_1__4 
       (.I0(\a6/k1a [2]),
        .I1(\a6/k4a [2]),
        .O(k5b[66]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[66]_i_1__5 
       (.I0(\a7/k1a [2]),
        .I1(\a7/k4a [2]),
        .O(k6b[66]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[66]_i_1__6 
       (.I0(\a8/k1a [2]),
        .I1(\a8/k4a [2]),
        .O(k7b[66]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[66]_i_1__7 
       (.I0(\a9/k1a [2]),
        .I1(\a9/k4a [2]),
        .O(k8b[66]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[67]_i_1 
       (.I0(\a1/k1a [3]),
        .I1(\a1/k4a [3]),
        .O(k0b[67]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[67]_i_1__0 
       (.I0(\a2/k1a [3]),
        .I1(\a2/k4a [3]),
        .O(k1b[67]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[67]_i_1__1 
       (.I0(\a3/k1a [3]),
        .I1(\a3/k4a [3]),
        .O(k2b[67]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[67]_i_1__2 
       (.I0(\a4/k1a [3]),
        .I1(\a4/k4a [3]),
        .O(k3b[67]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[67]_i_1__3 
       (.I0(\a5/k1a [3]),
        .I1(\a5/k4a [3]),
        .O(k4b[67]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[67]_i_1__4 
       (.I0(\a6/k1a [3]),
        .I1(\a6/k4a [3]),
        .O(k5b[67]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[67]_i_1__5 
       (.I0(\a7/k1a [3]),
        .I1(\a7/k4a [3]),
        .O(k6b[67]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[67]_i_1__6 
       (.I0(\a8/k1a [3]),
        .I1(\a8/k4a [3]),
        .O(k7b[67]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[67]_i_1__7 
       (.I0(\a9/k1a [3]),
        .I1(\a9/k4a [3]),
        .O(k8b[67]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[68]_i_1 
       (.I0(\a1/k1a [4]),
        .I1(\a1/k4a [4]),
        .O(k0b[68]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[68]_i_1__0 
       (.I0(\a2/k1a [4]),
        .I1(\a2/k4a [4]),
        .O(k1b[68]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[68]_i_1__1 
       (.I0(\a3/k1a [4]),
        .I1(\a3/k4a [4]),
        .O(k2b[68]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[68]_i_1__2 
       (.I0(\a4/k1a [4]),
        .I1(\a4/k4a [4]),
        .O(k3b[68]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[68]_i_1__3 
       (.I0(\a5/k1a [4]),
        .I1(\a5/k4a [4]),
        .O(k4b[68]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[68]_i_1__4 
       (.I0(\a6/k1a [4]),
        .I1(\a6/k4a [4]),
        .O(k5b[68]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[68]_i_1__5 
       (.I0(\a7/k1a [4]),
        .I1(\a7/k4a [4]),
        .O(k6b[68]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[68]_i_1__6 
       (.I0(\a8/k1a [4]),
        .I1(\a8/k4a [4]),
        .O(k7b[68]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[68]_i_1__7 
       (.I0(\a9/k1a [4]),
        .I1(\a9/k4a [4]),
        .O(k8b[68]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[69]_i_1 
       (.I0(\a1/k1a [5]),
        .I1(\a1/k4a [5]),
        .O(k0b[69]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[69]_i_1__0 
       (.I0(\a2/k1a [5]),
        .I1(\a2/k4a [5]),
        .O(k1b[69]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[69]_i_1__1 
       (.I0(\a3/k1a [5]),
        .I1(\a3/k4a [5]),
        .O(k2b[69]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[69]_i_1__2 
       (.I0(\a4/k1a [5]),
        .I1(\a4/k4a [5]),
        .O(k3b[69]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[69]_i_1__3 
       (.I0(\a5/k1a [5]),
        .I1(\a5/k4a [5]),
        .O(k4b[69]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[69]_i_1__4 
       (.I0(\a6/k1a [5]),
        .I1(\a6/k4a [5]),
        .O(k5b[69]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[69]_i_1__5 
       (.I0(\a7/k1a [5]),
        .I1(\a7/k4a [5]),
        .O(k6b[69]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[69]_i_1__6 
       (.I0(\a8/k1a [5]),
        .I1(\a8/k4a [5]),
        .O(k7b[69]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[69]_i_1__7 
       (.I0(\a9/k1a [5]),
        .I1(\a9/k4a [5]),
        .O(k8b[69]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[6]_i_1 
       (.I0(\a1/k3a [6]),
        .I1(\a1/k4a [6]),
        .O(k0b[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[6]_i_1__0 
       (.I0(\a2/k3a [6]),
        .I1(\a2/k4a [6]),
        .O(k1b[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[6]_i_1__1 
       (.I0(\a3/k3a [6]),
        .I1(\a3/k4a [6]),
        .O(k2b[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[6]_i_1__2 
       (.I0(\a4/k3a [6]),
        .I1(\a4/k4a [6]),
        .O(k3b[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[6]_i_1__3 
       (.I0(\a5/k3a [6]),
        .I1(\a5/k4a [6]),
        .O(k4b[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[6]_i_1__4 
       (.I0(\a6/k3a [6]),
        .I1(\a6/k4a [6]),
        .O(k5b[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[6]_i_1__5 
       (.I0(\a7/k3a [6]),
        .I1(\a7/k4a [6]),
        .O(k6b[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[6]_i_1__6 
       (.I0(\a8/k3a [6]),
        .I1(\a8/k4a [6]),
        .O(k7b[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[6]_i_1__7 
       (.I0(\a9/k3a [6]),
        .I1(\a9/k4a [6]),
        .O(k8b[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[70]_i_1 
       (.I0(\a1/k1a [6]),
        .I1(\a1/k4a [6]),
        .O(k0b[70]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[70]_i_1__0 
       (.I0(\a2/k1a [6]),
        .I1(\a2/k4a [6]),
        .O(k1b[70]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[70]_i_1__1 
       (.I0(\a3/k1a [6]),
        .I1(\a3/k4a [6]),
        .O(k2b[70]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[70]_i_1__2 
       (.I0(\a4/k1a [6]),
        .I1(\a4/k4a [6]),
        .O(k3b[70]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[70]_i_1__3 
       (.I0(\a5/k1a [6]),
        .I1(\a5/k4a [6]),
        .O(k4b[70]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[70]_i_1__4 
       (.I0(\a6/k1a [6]),
        .I1(\a6/k4a [6]),
        .O(k5b[70]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[70]_i_1__5 
       (.I0(\a7/k1a [6]),
        .I1(\a7/k4a [6]),
        .O(k6b[70]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[70]_i_1__6 
       (.I0(\a8/k1a [6]),
        .I1(\a8/k4a [6]),
        .O(k7b[70]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[70]_i_1__7 
       (.I0(\a9/k1a [6]),
        .I1(\a9/k4a [6]),
        .O(k8b[70]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[71]_i_1 
       (.I0(\a1/k1a [7]),
        .I1(\a1/k4a [7]),
        .O(k0b[71]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[71]_i_1__0 
       (.I0(\a2/k1a [7]),
        .I1(\a2/k4a [7]),
        .O(k1b[71]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[71]_i_1__1 
       (.I0(\a3/k1a [7]),
        .I1(\a3/k4a [7]),
        .O(k2b[71]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[71]_i_1__2 
       (.I0(\a4/k1a [7]),
        .I1(\a4/k4a [7]),
        .O(k3b[71]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[71]_i_1__3 
       (.I0(\a5/k1a [7]),
        .I1(\a5/k4a [7]),
        .O(k4b[71]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[71]_i_1__4 
       (.I0(\a6/k1a [7]),
        .I1(\a6/k4a [7]),
        .O(k5b[71]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[71]_i_1__5 
       (.I0(\a7/k1a [7]),
        .I1(\a7/k4a [7]),
        .O(k6b[71]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[71]_i_1__6 
       (.I0(\a8/k1a [7]),
        .I1(\a8/k4a [7]),
        .O(k7b[71]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[71]_i_1__7 
       (.I0(\a9/k1a [7]),
        .I1(\a9/k4a [7]),
        .O(k8b[71]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[72]_i_1 
       (.I0(\a1/k1a [8]),
        .I1(\a1/k4a [8]),
        .O(k0b[72]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[72]_i_1__0 
       (.I0(\a2/k1a [8]),
        .I1(\a2/k4a [8]),
        .O(k1b[72]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[72]_i_1__1 
       (.I0(\a3/k1a [8]),
        .I1(\a3/k4a [8]),
        .O(k2b[72]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[72]_i_1__2 
       (.I0(\a4/k1a [8]),
        .I1(\a4/k4a [8]),
        .O(k3b[72]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[72]_i_1__3 
       (.I0(\a5/k1a [8]),
        .I1(\a5/k4a [8]),
        .O(k4b[72]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[72]_i_1__4 
       (.I0(\a6/k1a [8]),
        .I1(\a6/k4a [8]),
        .O(k5b[72]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[72]_i_1__5 
       (.I0(\a7/k1a [8]),
        .I1(\a7/k4a [8]),
        .O(k6b[72]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[72]_i_1__6 
       (.I0(\a8/k1a [8]),
        .I1(\a8/k4a [8]),
        .O(k7b[72]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[72]_i_1__7 
       (.I0(\a9/k1a [8]),
        .I1(\a9/k4a [8]),
        .O(k8b[72]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[73]_i_1 
       (.I0(\a1/k1a [9]),
        .I1(\a1/k4a [9]),
        .O(k0b[73]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[73]_i_1__0 
       (.I0(\a2/k1a [9]),
        .I1(\a2/k4a [9]),
        .O(k1b[73]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[73]_i_1__1 
       (.I0(\a3/k1a [9]),
        .I1(\a3/k4a [9]),
        .O(k2b[73]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[73]_i_1__2 
       (.I0(\a4/k1a [9]),
        .I1(\a4/k4a [9]),
        .O(k3b[73]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[73]_i_1__3 
       (.I0(\a5/k1a [9]),
        .I1(\a5/k4a [9]),
        .O(k4b[73]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[73]_i_1__4 
       (.I0(\a6/k1a [9]),
        .I1(\a6/k4a [9]),
        .O(k5b[73]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[73]_i_1__5 
       (.I0(\a7/k1a [9]),
        .I1(\a7/k4a [9]),
        .O(k6b[73]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[73]_i_1__6 
       (.I0(\a8/k1a [9]),
        .I1(\a8/k4a [9]),
        .O(k7b[73]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[73]_i_1__7 
       (.I0(\a9/k1a [9]),
        .I1(\a9/k4a [9]),
        .O(k8b[73]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[74]_i_1 
       (.I0(\a1/k1a [10]),
        .I1(\a1/k4a [10]),
        .O(k0b[74]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[74]_i_1__0 
       (.I0(\a2/k1a [10]),
        .I1(\a2/k4a [10]),
        .O(k1b[74]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[74]_i_1__1 
       (.I0(\a3/k1a [10]),
        .I1(\a3/k4a [10]),
        .O(k2b[74]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[74]_i_1__2 
       (.I0(\a4/k1a [10]),
        .I1(\a4/k4a [10]),
        .O(k3b[74]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[74]_i_1__3 
       (.I0(\a5/k1a [10]),
        .I1(\a5/k4a [10]),
        .O(k4b[74]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[74]_i_1__4 
       (.I0(\a6/k1a [10]),
        .I1(\a6/k4a [10]),
        .O(k5b[74]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[74]_i_1__5 
       (.I0(\a7/k1a [10]),
        .I1(\a7/k4a [10]),
        .O(k6b[74]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[74]_i_1__6 
       (.I0(\a8/k1a [10]),
        .I1(\a8/k4a [10]),
        .O(k7b[74]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[74]_i_1__7 
       (.I0(\a9/k1a [10]),
        .I1(\a9/k4a [10]),
        .O(k8b[74]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[75]_i_1 
       (.I0(\a1/k1a [11]),
        .I1(\a1/k4a [11]),
        .O(k0b[75]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[75]_i_1__0 
       (.I0(\a2/k1a [11]),
        .I1(\a2/k4a [11]),
        .O(k1b[75]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[75]_i_1__1 
       (.I0(\a3/k1a [11]),
        .I1(\a3/k4a [11]),
        .O(k2b[75]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[75]_i_1__2 
       (.I0(\a4/k1a [11]),
        .I1(\a4/k4a [11]),
        .O(k3b[75]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[75]_i_1__3 
       (.I0(\a5/k1a [11]),
        .I1(\a5/k4a [11]),
        .O(k4b[75]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[75]_i_1__4 
       (.I0(\a6/k1a [11]),
        .I1(\a6/k4a [11]),
        .O(k5b[75]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[75]_i_1__5 
       (.I0(\a7/k1a [11]),
        .I1(\a7/k4a [11]),
        .O(k6b[75]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[75]_i_1__6 
       (.I0(\a8/k1a [11]),
        .I1(\a8/k4a [11]),
        .O(k7b[75]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[75]_i_1__7 
       (.I0(\a9/k1a [11]),
        .I1(\a9/k4a [11]),
        .O(k8b[75]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[76]_i_1 
       (.I0(\a1/k1a [12]),
        .I1(\a1/k4a [12]),
        .O(k0b[76]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[76]_i_1__0 
       (.I0(\a2/k1a [12]),
        .I1(\a2/k4a [12]),
        .O(k1b[76]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[76]_i_1__1 
       (.I0(\a3/k1a [12]),
        .I1(\a3/k4a [12]),
        .O(k2b[76]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[76]_i_1__2 
       (.I0(\a4/k1a [12]),
        .I1(\a4/k4a [12]),
        .O(k3b[76]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[76]_i_1__3 
       (.I0(\a5/k1a [12]),
        .I1(\a5/k4a [12]),
        .O(k4b[76]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[76]_i_1__4 
       (.I0(\a6/k1a [12]),
        .I1(\a6/k4a [12]),
        .O(k5b[76]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[76]_i_1__5 
       (.I0(\a7/k1a [12]),
        .I1(\a7/k4a [12]),
        .O(k6b[76]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[76]_i_1__6 
       (.I0(\a8/k1a [12]),
        .I1(\a8/k4a [12]),
        .O(k7b[76]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[76]_i_1__7 
       (.I0(\a9/k1a [12]),
        .I1(\a9/k4a [12]),
        .O(k8b[76]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[77]_i_1 
       (.I0(\a1/k1a [13]),
        .I1(\a1/k4a [13]),
        .O(k0b[77]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[77]_i_1__0 
       (.I0(\a2/k1a [13]),
        .I1(\a2/k4a [13]),
        .O(k1b[77]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[77]_i_1__1 
       (.I0(\a3/k1a [13]),
        .I1(\a3/k4a [13]),
        .O(k2b[77]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[77]_i_1__2 
       (.I0(\a4/k1a [13]),
        .I1(\a4/k4a [13]),
        .O(k3b[77]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[77]_i_1__3 
       (.I0(\a5/k1a [13]),
        .I1(\a5/k4a [13]),
        .O(k4b[77]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[77]_i_1__4 
       (.I0(\a6/k1a [13]),
        .I1(\a6/k4a [13]),
        .O(k5b[77]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[77]_i_1__5 
       (.I0(\a7/k1a [13]),
        .I1(\a7/k4a [13]),
        .O(k6b[77]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[77]_i_1__6 
       (.I0(\a8/k1a [13]),
        .I1(\a8/k4a [13]),
        .O(k7b[77]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[77]_i_1__7 
       (.I0(\a9/k1a [13]),
        .I1(\a9/k4a [13]),
        .O(k8b[77]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[78]_i_1 
       (.I0(\a1/k1a [14]),
        .I1(\a1/k4a [14]),
        .O(k0b[78]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[78]_i_1__0 
       (.I0(\a2/k1a [14]),
        .I1(\a2/k4a [14]),
        .O(k1b[78]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[78]_i_1__1 
       (.I0(\a3/k1a [14]),
        .I1(\a3/k4a [14]),
        .O(k2b[78]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[78]_i_1__2 
       (.I0(\a4/k1a [14]),
        .I1(\a4/k4a [14]),
        .O(k3b[78]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[78]_i_1__3 
       (.I0(\a5/k1a [14]),
        .I1(\a5/k4a [14]),
        .O(k4b[78]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[78]_i_1__4 
       (.I0(\a6/k1a [14]),
        .I1(\a6/k4a [14]),
        .O(k5b[78]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[78]_i_1__5 
       (.I0(\a7/k1a [14]),
        .I1(\a7/k4a [14]),
        .O(k6b[78]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[78]_i_1__6 
       (.I0(\a8/k1a [14]),
        .I1(\a8/k4a [14]),
        .O(k7b[78]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[78]_i_1__7 
       (.I0(\a9/k1a [14]),
        .I1(\a9/k4a [14]),
        .O(k8b[78]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[79]_i_1 
       (.I0(\a1/k1a [15]),
        .I1(\a1/k4a [15]),
        .O(k0b[79]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[79]_i_1__0 
       (.I0(\a2/k1a [15]),
        .I1(\a2/k4a [15]),
        .O(k1b[79]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[79]_i_1__1 
       (.I0(\a3/k1a [15]),
        .I1(\a3/k4a [15]),
        .O(k2b[79]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[79]_i_1__2 
       (.I0(\a4/k1a [15]),
        .I1(\a4/k4a [15]),
        .O(k3b[79]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[79]_i_1__3 
       (.I0(\a5/k1a [15]),
        .I1(\a5/k4a [15]),
        .O(k4b[79]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[79]_i_1__4 
       (.I0(\a6/k1a [15]),
        .I1(\a6/k4a [15]),
        .O(k5b[79]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[79]_i_1__5 
       (.I0(\a7/k1a [15]),
        .I1(\a7/k4a [15]),
        .O(k6b[79]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[79]_i_1__6 
       (.I0(\a8/k1a [15]),
        .I1(\a8/k4a [15]),
        .O(k7b[79]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[79]_i_1__7 
       (.I0(\a9/k1a [15]),
        .I1(\a9/k4a [15]),
        .O(k8b[79]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[7]_i_1 
       (.I0(\a1/k3a [7]),
        .I1(\a1/k4a [7]),
        .O(k0b[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[7]_i_1__0 
       (.I0(\a2/k3a [7]),
        .I1(\a2/k4a [7]),
        .O(k1b[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[7]_i_1__1 
       (.I0(\a3/k3a [7]),
        .I1(\a3/k4a [7]),
        .O(k2b[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[7]_i_1__2 
       (.I0(\a4/k3a [7]),
        .I1(\a4/k4a [7]),
        .O(k3b[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[7]_i_1__3 
       (.I0(\a5/k3a [7]),
        .I1(\a5/k4a [7]),
        .O(k4b[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[7]_i_1__4 
       (.I0(\a6/k3a [7]),
        .I1(\a6/k4a [7]),
        .O(k5b[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[7]_i_1__5 
       (.I0(\a7/k3a [7]),
        .I1(\a7/k4a [7]),
        .O(k6b[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[7]_i_1__6 
       (.I0(\a8/k3a [7]),
        .I1(\a8/k4a [7]),
        .O(k7b[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[7]_i_1__7 
       (.I0(\a9/k3a [7]),
        .I1(\a9/k4a [7]),
        .O(k8b[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[80]_i_1 
       (.I0(\a1/k1a [16]),
        .I1(\a1/k4a [16]),
        .O(k0b[80]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[80]_i_1__0 
       (.I0(\a2/k1a [16]),
        .I1(\a2/k4a [16]),
        .O(k1b[80]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[80]_i_1__1 
       (.I0(\a3/k1a [16]),
        .I1(\a3/k4a [16]),
        .O(k2b[80]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[80]_i_1__2 
       (.I0(\a4/k1a [16]),
        .I1(\a4/k4a [16]),
        .O(k3b[80]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[80]_i_1__3 
       (.I0(\a5/k1a [16]),
        .I1(\a5/k4a [16]),
        .O(k4b[80]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[80]_i_1__4 
       (.I0(\a6/k1a [16]),
        .I1(\a6/k4a [16]),
        .O(k5b[80]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[80]_i_1__5 
       (.I0(\a7/k1a [16]),
        .I1(\a7/k4a [16]),
        .O(k6b[80]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[80]_i_1__6 
       (.I0(\a8/k1a [16]),
        .I1(\a8/k4a [16]),
        .O(k7b[80]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[80]_i_1__7 
       (.I0(\a9/k1a [16]),
        .I1(\a9/k4a [16]),
        .O(k8b[80]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[81]_i_1 
       (.I0(\a1/k1a [17]),
        .I1(\a1/k4a [17]),
        .O(k0b[81]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[81]_i_1__0 
       (.I0(\a2/k1a [17]),
        .I1(\a2/k4a [17]),
        .O(k1b[81]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[81]_i_1__1 
       (.I0(\a3/k1a [17]),
        .I1(\a3/k4a [17]),
        .O(k2b[81]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[81]_i_1__2 
       (.I0(\a4/k1a [17]),
        .I1(\a4/k4a [17]),
        .O(k3b[81]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[81]_i_1__3 
       (.I0(\a5/k1a [17]),
        .I1(\a5/k4a [17]),
        .O(k4b[81]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[81]_i_1__4 
       (.I0(\a6/k1a [17]),
        .I1(\a6/k4a [17]),
        .O(k5b[81]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[81]_i_1__5 
       (.I0(\a7/k1a [17]),
        .I1(\a7/k4a [17]),
        .O(k6b[81]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[81]_i_1__6 
       (.I0(\a8/k1a [17]),
        .I1(\a8/k4a [17]),
        .O(k7b[81]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[81]_i_1__7 
       (.I0(\a9/k1a [17]),
        .I1(\a9/k4a [17]),
        .O(k8b[81]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[82]_i_1 
       (.I0(\a1/k1a [18]),
        .I1(\a1/k4a [18]),
        .O(k0b[82]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[82]_i_1__0 
       (.I0(\a2/k1a [18]),
        .I1(\a2/k4a [18]),
        .O(k1b[82]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[82]_i_1__1 
       (.I0(\a3/k1a [18]),
        .I1(\a3/k4a [18]),
        .O(k2b[82]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[82]_i_1__2 
       (.I0(\a4/k1a [18]),
        .I1(\a4/k4a [18]),
        .O(k3b[82]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[82]_i_1__3 
       (.I0(\a5/k1a [18]),
        .I1(\a5/k4a [18]),
        .O(k4b[82]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[82]_i_1__4 
       (.I0(\a6/k1a [18]),
        .I1(\a6/k4a [18]),
        .O(k5b[82]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[82]_i_1__5 
       (.I0(\a7/k1a [18]),
        .I1(\a7/k4a [18]),
        .O(k6b[82]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[82]_i_1__6 
       (.I0(\a8/k1a [18]),
        .I1(\a8/k4a [18]),
        .O(k7b[82]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[82]_i_1__7 
       (.I0(\a9/k1a [18]),
        .I1(\a9/k4a [18]),
        .O(k8b[82]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[83]_i_1 
       (.I0(\a1/k1a [19]),
        .I1(\a1/k4a [19]),
        .O(k0b[83]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[83]_i_1__0 
       (.I0(\a2/k1a [19]),
        .I1(\a2/k4a [19]),
        .O(k1b[83]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[83]_i_1__1 
       (.I0(\a3/k1a [19]),
        .I1(\a3/k4a [19]),
        .O(k2b[83]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[83]_i_1__2 
       (.I0(\a4/k1a [19]),
        .I1(\a4/k4a [19]),
        .O(k3b[83]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[83]_i_1__3 
       (.I0(\a5/k1a [19]),
        .I1(\a5/k4a [19]),
        .O(k4b[83]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[83]_i_1__4 
       (.I0(\a6/k1a [19]),
        .I1(\a6/k4a [19]),
        .O(k5b[83]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[83]_i_1__5 
       (.I0(\a7/k1a [19]),
        .I1(\a7/k4a [19]),
        .O(k6b[83]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[83]_i_1__6 
       (.I0(\a8/k1a [19]),
        .I1(\a8/k4a [19]),
        .O(k7b[83]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[83]_i_1__7 
       (.I0(\a9/k1a [19]),
        .I1(\a9/k4a [19]),
        .O(k8b[83]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[84]_i_1 
       (.I0(\a1/k1a [20]),
        .I1(\a1/k4a [20]),
        .O(k0b[84]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[84]_i_1__0 
       (.I0(\a2/k1a [20]),
        .I1(\a2/k4a [20]),
        .O(k1b[84]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[84]_i_1__1 
       (.I0(\a3/k1a [20]),
        .I1(\a3/k4a [20]),
        .O(k2b[84]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[84]_i_1__2 
       (.I0(\a4/k1a [20]),
        .I1(\a4/k4a [20]),
        .O(k3b[84]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[84]_i_1__3 
       (.I0(\a5/k1a [20]),
        .I1(\a5/k4a [20]),
        .O(k4b[84]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[84]_i_1__4 
       (.I0(\a6/k1a [20]),
        .I1(\a6/k4a [20]),
        .O(k5b[84]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[84]_i_1__5 
       (.I0(\a7/k1a [20]),
        .I1(\a7/k4a [20]),
        .O(k6b[84]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[84]_i_1__6 
       (.I0(\a8/k1a [20]),
        .I1(\a8/k4a [20]),
        .O(k7b[84]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[84]_i_1__7 
       (.I0(\a9/k1a [20]),
        .I1(\a9/k4a [20]),
        .O(k8b[84]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[85]_i_1 
       (.I0(\a1/k1a [21]),
        .I1(\a1/k4a [21]),
        .O(k0b[85]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[85]_i_1__0 
       (.I0(\a2/k1a [21]),
        .I1(\a2/k4a [21]),
        .O(k1b[85]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[85]_i_1__1 
       (.I0(\a3/k1a [21]),
        .I1(\a3/k4a [21]),
        .O(k2b[85]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[85]_i_1__2 
       (.I0(\a4/k1a [21]),
        .I1(\a4/k4a [21]),
        .O(k3b[85]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[85]_i_1__3 
       (.I0(\a5/k1a [21]),
        .I1(\a5/k4a [21]),
        .O(k4b[85]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[85]_i_1__4 
       (.I0(\a6/k1a [21]),
        .I1(\a6/k4a [21]),
        .O(k5b[85]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[85]_i_1__5 
       (.I0(\a7/k1a [21]),
        .I1(\a7/k4a [21]),
        .O(k6b[85]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[85]_i_1__6 
       (.I0(\a8/k1a [21]),
        .I1(\a8/k4a [21]),
        .O(k7b[85]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[85]_i_1__7 
       (.I0(\a9/k1a [21]),
        .I1(\a9/k4a [21]),
        .O(k8b[85]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[86]_i_1 
       (.I0(\a1/k1a [22]),
        .I1(\a1/k4a [22]),
        .O(k0b[86]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[86]_i_1__0 
       (.I0(\a2/k1a [22]),
        .I1(\a2/k4a [22]),
        .O(k1b[86]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[86]_i_1__1 
       (.I0(\a3/k1a [22]),
        .I1(\a3/k4a [22]),
        .O(k2b[86]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[86]_i_1__2 
       (.I0(\a4/k1a [22]),
        .I1(\a4/k4a [22]),
        .O(k3b[86]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[86]_i_1__3 
       (.I0(\a5/k1a [22]),
        .I1(\a5/k4a [22]),
        .O(k4b[86]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[86]_i_1__4 
       (.I0(\a6/k1a [22]),
        .I1(\a6/k4a [22]),
        .O(k5b[86]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[86]_i_1__5 
       (.I0(\a7/k1a [22]),
        .I1(\a7/k4a [22]),
        .O(k6b[86]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[86]_i_1__6 
       (.I0(\a8/k1a [22]),
        .I1(\a8/k4a [22]),
        .O(k7b[86]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[86]_i_1__7 
       (.I0(\a9/k1a [22]),
        .I1(\a9/k4a [22]),
        .O(k8b[86]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[87]_i_1 
       (.I0(\a1/k1a [23]),
        .I1(\a1/k4a [23]),
        .O(k0b[87]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[87]_i_1__0 
       (.I0(\a2/k1a [23]),
        .I1(\a2/k4a [23]),
        .O(k1b[87]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[87]_i_1__1 
       (.I0(\a3/k1a [23]),
        .I1(\a3/k4a [23]),
        .O(k2b[87]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[87]_i_1__2 
       (.I0(\a4/k1a [23]),
        .I1(\a4/k4a [23]),
        .O(k3b[87]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[87]_i_1__3 
       (.I0(\a5/k1a [23]),
        .I1(\a5/k4a [23]),
        .O(k4b[87]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[87]_i_1__4 
       (.I0(\a6/k1a [23]),
        .I1(\a6/k4a [23]),
        .O(k5b[87]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[87]_i_1__5 
       (.I0(\a7/k1a [23]),
        .I1(\a7/k4a [23]),
        .O(k6b[87]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[87]_i_1__6 
       (.I0(\a8/k1a [23]),
        .I1(\a8/k4a [23]),
        .O(k7b[87]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[87]_i_1__7 
       (.I0(\a9/k1a [23]),
        .I1(\a9/k4a [23]),
        .O(k8b[87]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[88]_i_1 
       (.I0(\a1/k1a [24]),
        .I1(\a1/k4a [24]),
        .O(k0b[88]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[88]_i_1__0 
       (.I0(\a2/k1a [24]),
        .I1(\a2/k4a [24]),
        .O(k1b[88]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[88]_i_1__1 
       (.I0(\a3/k1a [24]),
        .I1(\a3/k4a [24]),
        .O(k2b[88]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[88]_i_1__2 
       (.I0(\a4/k1a [24]),
        .I1(\a4/k4a [24]),
        .O(k3b[88]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[88]_i_1__3 
       (.I0(\a5/k1a [24]),
        .I1(\a5/k4a [24]),
        .O(k4b[88]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[88]_i_1__4 
       (.I0(\a6/k1a [24]),
        .I1(\a6/k4a [24]),
        .O(k5b[88]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[88]_i_1__5 
       (.I0(\a7/k1a [24]),
        .I1(\a7/k4a [24]),
        .O(k6b[88]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[88]_i_1__6 
       (.I0(\a8/k1a [24]),
        .I1(\a8/k4a [24]),
        .O(k7b[88]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[88]_i_1__7 
       (.I0(\a9/k1a [24]),
        .I1(\a9/k4a [24]),
        .O(k8b[88]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[89]_i_1 
       (.I0(\a1/k1a [25]),
        .I1(\a1/k4a [25]),
        .O(k0b[89]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[89]_i_1__0 
       (.I0(\a2/k1a [25]),
        .I1(\a2/k4a [25]),
        .O(k1b[89]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[89]_i_1__1 
       (.I0(\a3/k1a [25]),
        .I1(\a3/k4a [25]),
        .O(k2b[89]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[89]_i_1__2 
       (.I0(\a4/k1a [25]),
        .I1(\a4/k4a [25]),
        .O(k3b[89]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[89]_i_1__3 
       (.I0(\a5/k1a [25]),
        .I1(\a5/k4a [25]),
        .O(k4b[89]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[89]_i_1__4 
       (.I0(\a6/k1a [25]),
        .I1(\a6/k4a [25]),
        .O(k5b[89]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[89]_i_1__5 
       (.I0(\a7/k1a [25]),
        .I1(\a7/k4a [25]),
        .O(k6b[89]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[89]_i_1__6 
       (.I0(\a8/k1a [25]),
        .I1(\a8/k4a [25]),
        .O(k7b[89]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[89]_i_1__7 
       (.I0(\a9/k1a [25]),
        .I1(\a9/k4a [25]),
        .O(k8b[89]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[8]_i_1 
       (.I0(\a1/k3a [8]),
        .I1(\a1/k4a [8]),
        .O(k0b[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[8]_i_1__0 
       (.I0(\a2/k3a [8]),
        .I1(\a2/k4a [8]),
        .O(k1b[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[8]_i_1__1 
       (.I0(\a3/k3a [8]),
        .I1(\a3/k4a [8]),
        .O(k2b[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[8]_i_1__2 
       (.I0(\a4/k3a [8]),
        .I1(\a4/k4a [8]),
        .O(k3b[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[8]_i_1__3 
       (.I0(\a5/k3a [8]),
        .I1(\a5/k4a [8]),
        .O(k4b[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[8]_i_1__4 
       (.I0(\a6/k3a [8]),
        .I1(\a6/k4a [8]),
        .O(k5b[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[8]_i_1__5 
       (.I0(\a7/k3a [8]),
        .I1(\a7/k4a [8]),
        .O(k6b[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[8]_i_1__6 
       (.I0(\a8/k3a [8]),
        .I1(\a8/k4a [8]),
        .O(k7b[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[8]_i_1__7 
       (.I0(\a9/k3a [8]),
        .I1(\a9/k4a [8]),
        .O(k8b[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[90]_i_1 
       (.I0(\a1/k1a [26]),
        .I1(\a1/k4a [26]),
        .O(k0b[90]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[90]_i_1__0 
       (.I0(\a2/k1a [26]),
        .I1(\a2/k4a [26]),
        .O(k1b[90]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[90]_i_1__1 
       (.I0(\a3/k1a [26]),
        .I1(\a3/k4a [26]),
        .O(k2b[90]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[90]_i_1__2 
       (.I0(\a4/k1a [26]),
        .I1(\a4/k4a [26]),
        .O(k3b[90]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[90]_i_1__3 
       (.I0(\a5/k1a [26]),
        .I1(\a5/k4a [26]),
        .O(k4b[90]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[90]_i_1__4 
       (.I0(\a6/k1a [26]),
        .I1(\a6/k4a [26]),
        .O(k5b[90]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[90]_i_1__5 
       (.I0(\a7/k1a [26]),
        .I1(\a7/k4a [26]),
        .O(k6b[90]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[90]_i_1__6 
       (.I0(\a8/k1a [26]),
        .I1(\a8/k4a [26]),
        .O(k7b[90]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[90]_i_1__7 
       (.I0(\a9/k1a [26]),
        .I1(\a9/k4a [26]),
        .O(k8b[90]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[91]_i_1 
       (.I0(\a1/k1a [27]),
        .I1(\a1/k4a [27]),
        .O(k0b[91]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[91]_i_1__0 
       (.I0(\a2/k1a [27]),
        .I1(\a2/k4a [27]),
        .O(k1b[91]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[91]_i_1__1 
       (.I0(\a3/k1a [27]),
        .I1(\a3/k4a [27]),
        .O(k2b[91]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[91]_i_1__2 
       (.I0(\a4/k1a [27]),
        .I1(\a4/k4a [27]),
        .O(k3b[91]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[91]_i_1__3 
       (.I0(\a5/k1a [27]),
        .I1(\a5/k4a [27]),
        .O(k4b[91]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[91]_i_1__4 
       (.I0(\a6/k1a [27]),
        .I1(\a6/k4a [27]),
        .O(k5b[91]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[91]_i_1__5 
       (.I0(\a7/k1a [27]),
        .I1(\a7/k4a [27]),
        .O(k6b[91]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[91]_i_1__6 
       (.I0(\a8/k1a [27]),
        .I1(\a8/k4a [27]),
        .O(k7b[91]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[91]_i_1__7 
       (.I0(\a9/k1a [27]),
        .I1(\a9/k4a [27]),
        .O(k8b[91]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[92]_i_1 
       (.I0(\a1/k1a [28]),
        .I1(\a1/k4a [28]),
        .O(k0b[92]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[92]_i_1__0 
       (.I0(\a2/k1a [28]),
        .I1(\a2/k4a [28]),
        .O(k1b[92]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[92]_i_1__1 
       (.I0(\a3/k1a [28]),
        .I1(\a3/k4a [28]),
        .O(k2b[92]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[92]_i_1__2 
       (.I0(\a4/k1a [28]),
        .I1(\a4/k4a [28]),
        .O(k3b[92]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[92]_i_1__3 
       (.I0(\a5/k1a [28]),
        .I1(\a5/k4a [28]),
        .O(k4b[92]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[92]_i_1__4 
       (.I0(\a6/k1a [28]),
        .I1(\a6/k4a [28]),
        .O(k5b[92]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[92]_i_1__5 
       (.I0(\a7/k1a [28]),
        .I1(\a7/k4a [28]),
        .O(k6b[92]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[92]_i_1__6 
       (.I0(\a8/k1a [28]),
        .I1(\a8/k4a [28]),
        .O(k7b[92]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[92]_i_1__7 
       (.I0(\a9/k1a [28]),
        .I1(\a9/k4a [28]),
        .O(k8b[92]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[93]_i_1 
       (.I0(\a1/k1a [29]),
        .I1(\a1/k4a [29]),
        .O(k0b[93]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[93]_i_1__0 
       (.I0(\a2/k1a [29]),
        .I1(\a2/k4a [29]),
        .O(k1b[93]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[93]_i_1__1 
       (.I0(\a3/k1a [29]),
        .I1(\a3/k4a [29]),
        .O(k2b[93]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[93]_i_1__2 
       (.I0(\a4/k1a [29]),
        .I1(\a4/k4a [29]),
        .O(k3b[93]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[93]_i_1__3 
       (.I0(\a5/k1a [29]),
        .I1(\a5/k4a [29]),
        .O(k4b[93]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[93]_i_1__4 
       (.I0(\a6/k1a [29]),
        .I1(\a6/k4a [29]),
        .O(k5b[93]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[93]_i_1__5 
       (.I0(\a7/k1a [29]),
        .I1(\a7/k4a [29]),
        .O(k6b[93]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[93]_i_1__6 
       (.I0(\a8/k1a [29]),
        .I1(\a8/k4a [29]),
        .O(k7b[93]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[93]_i_1__7 
       (.I0(\a9/k1a [29]),
        .I1(\a9/k4a [29]),
        .O(k8b[93]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[94]_i_1 
       (.I0(\a1/k1a [30]),
        .I1(\a1/k4a [30]),
        .O(k0b[94]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[94]_i_1__0 
       (.I0(\a2/k1a [30]),
        .I1(\a2/k4a [30]),
        .O(k1b[94]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[94]_i_1__1 
       (.I0(\a3/k1a [30]),
        .I1(\a3/k4a [30]),
        .O(k2b[94]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[94]_i_1__2 
       (.I0(\a4/k1a [30]),
        .I1(\a4/k4a [30]),
        .O(k3b[94]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[94]_i_1__3 
       (.I0(\a5/k1a [30]),
        .I1(\a5/k4a [30]),
        .O(k4b[94]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[94]_i_1__4 
       (.I0(\a6/k1a [30]),
        .I1(\a6/k4a [30]),
        .O(k5b[94]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[94]_i_1__5 
       (.I0(\a7/k1a [30]),
        .I1(\a7/k4a [30]),
        .O(k6b[94]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[94]_i_1__6 
       (.I0(\a8/k1a [30]),
        .I1(\a8/k4a [30]),
        .O(k7b[94]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[94]_i_1__7 
       (.I0(\a9/k1a [30]),
        .I1(\a9/k4a [30]),
        .O(k8b[94]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[95]_i_1 
       (.I0(\a1/k1a [31]),
        .I1(\a1/k4a [31]),
        .O(k0b[95]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[95]_i_1__0 
       (.I0(\a2/k1a [31]),
        .I1(\a2/k4a [31]),
        .O(k1b[95]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[95]_i_1__1 
       (.I0(\a3/k1a [31]),
        .I1(\a3/k4a [31]),
        .O(k2b[95]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[95]_i_1__2 
       (.I0(\a4/k1a [31]),
        .I1(\a4/k4a [31]),
        .O(k3b[95]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[95]_i_1__3 
       (.I0(\a5/k1a [31]),
        .I1(\a5/k4a [31]),
        .O(k4b[95]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[95]_i_1__4 
       (.I0(\a6/k1a [31]),
        .I1(\a6/k4a [31]),
        .O(k5b[95]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[95]_i_1__5 
       (.I0(\a7/k1a [31]),
        .I1(\a7/k4a [31]),
        .O(k6b[95]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[95]_i_1__6 
       (.I0(\a8/k1a [31]),
        .I1(\a8/k4a [31]),
        .O(k7b[95]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[95]_i_1__7 
       (.I0(\a9/k1a [31]),
        .I1(\a9/k4a [31]),
        .O(k8b[95]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[96]_i_1 
       (.I0(\a1/k0a [0]),
        .I1(\a1/k4a [0]),
        .O(k0b[96]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[96]_i_1__0 
       (.I0(\a2/k0a [0]),
        .I1(\a2/k4a [0]),
        .O(k1b[96]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[96]_i_1__1 
       (.I0(\a3/k0a [0]),
        .I1(\a3/k4a [0]),
        .O(k2b[96]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[96]_i_1__2 
       (.I0(\a4/k0a [0]),
        .I1(\a4/k4a [0]),
        .O(k3b[96]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[96]_i_1__3 
       (.I0(\a5/k0a [0]),
        .I1(\a5/k4a [0]),
        .O(k4b[96]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[96]_i_1__4 
       (.I0(\a6/k0a [0]),
        .I1(\a6/k4a [0]),
        .O(k5b[96]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[96]_i_1__5 
       (.I0(\a7/k0a [0]),
        .I1(\a7/k4a [0]),
        .O(k6b[96]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[96]_i_1__6 
       (.I0(\a8/k0a [0]),
        .I1(\a8/k4a [0]),
        .O(k7b[96]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[96]_i_1__7 
       (.I0(\a9/k0a [0]),
        .I1(\a9/k4a [0]),
        .O(k8b[96]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[97]_i_1 
       (.I0(\a1/k0a [1]),
        .I1(\a1/k4a [1]),
        .O(k0b[97]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[97]_i_1__0 
       (.I0(\a2/k0a [1]),
        .I1(\a2/k4a [1]),
        .O(k1b[97]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[97]_i_1__1 
       (.I0(\a3/k0a [1]),
        .I1(\a3/k4a [1]),
        .O(k2b[97]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[97]_i_1__2 
       (.I0(\a4/k0a [1]),
        .I1(\a4/k4a [1]),
        .O(k3b[97]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[97]_i_1__3 
       (.I0(\a5/k0a [1]),
        .I1(\a5/k4a [1]),
        .O(k4b[97]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[97]_i_1__4 
       (.I0(\a6/k0a [1]),
        .I1(\a6/k4a [1]),
        .O(k5b[97]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[97]_i_1__5 
       (.I0(\a7/k0a [1]),
        .I1(\a7/k4a [1]),
        .O(k6b[97]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[97]_i_1__6 
       (.I0(\a8/k0a [1]),
        .I1(\a8/k4a [1]),
        .O(k7b[97]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[97]_i_1__7 
       (.I0(\a9/k0a [1]),
        .I1(\a9/k4a [1]),
        .O(k8b[97]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[98]_i_1 
       (.I0(\a1/k0a [2]),
        .I1(\a1/k4a [2]),
        .O(k0b[98]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[98]_i_1__0 
       (.I0(\a2/k0a [2]),
        .I1(\a2/k4a [2]),
        .O(k1b[98]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[98]_i_1__1 
       (.I0(\a3/k0a [2]),
        .I1(\a3/k4a [2]),
        .O(k2b[98]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[98]_i_1__2 
       (.I0(\a4/k0a [2]),
        .I1(\a4/k4a [2]),
        .O(k3b[98]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[98]_i_1__3 
       (.I0(\a5/k0a [2]),
        .I1(\a5/k4a [2]),
        .O(k4b[98]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[98]_i_1__4 
       (.I0(\a6/k0a [2]),
        .I1(\a6/k4a [2]),
        .O(k5b[98]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[98]_i_1__5 
       (.I0(\a7/k0a [2]),
        .I1(\a7/k4a [2]),
        .O(k6b[98]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[98]_i_1__6 
       (.I0(\a8/k0a [2]),
        .I1(\a8/k4a [2]),
        .O(k7b[98]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[98]_i_1__7 
       (.I0(\a9/k0a [2]),
        .I1(\a9/k4a [2]),
        .O(k8b[98]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[99]_i_1 
       (.I0(\a1/k0a [3]),
        .I1(\a1/k4a [3]),
        .O(k0b[99]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[99]_i_1__0 
       (.I0(\a2/k0a [3]),
        .I1(\a2/k4a [3]),
        .O(k1b[99]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[99]_i_1__1 
       (.I0(\a3/k0a [3]),
        .I1(\a3/k4a [3]),
        .O(k2b[99]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[99]_i_1__2 
       (.I0(\a4/k0a [3]),
        .I1(\a4/k4a [3]),
        .O(k3b[99]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[99]_i_1__3 
       (.I0(\a5/k0a [3]),
        .I1(\a5/k4a [3]),
        .O(k4b[99]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[99]_i_1__4 
       (.I0(\a6/k0a [3]),
        .I1(\a6/k4a [3]),
        .O(k5b[99]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[99]_i_1__5 
       (.I0(\a7/k0a [3]),
        .I1(\a7/k4a [3]),
        .O(k6b[99]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[99]_i_1__6 
       (.I0(\a8/k0a [3]),
        .I1(\a8/k4a [3]),
        .O(k7b[99]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[99]_i_1__7 
       (.I0(\a9/k0a [3]),
        .I1(\a9/k4a [3]),
        .O(k8b[99]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[9]_i_1 
       (.I0(\a1/k3a [9]),
        .I1(\a1/k4a [9]),
        .O(k0b[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[9]_i_1__0 
       (.I0(\a2/k3a [9]),
        .I1(\a2/k4a [9]),
        .O(k1b[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[9]_i_1__1 
       (.I0(\a3/k3a [9]),
        .I1(\a3/k4a [9]),
        .O(k2b[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[9]_i_1__2 
       (.I0(\a4/k3a [9]),
        .I1(\a4/k4a [9]),
        .O(k3b[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[9]_i_1__3 
       (.I0(\a5/k3a [9]),
        .I1(\a5/k4a [9]),
        .O(k4b[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[9]_i_1__4 
       (.I0(\a6/k3a [9]),
        .I1(\a6/k4a [9]),
        .O(k5b[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[9]_i_1__5 
       (.I0(\a7/k3a [9]),
        .I1(\a7/k4a [9]),
        .O(k6b[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[9]_i_1__6 
       (.I0(\a8/k3a [9]),
        .I1(\a8/k4a [9]),
        .O(k7b[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \out_1[9]_i_1__7 
       (.I0(\a9/k3a [9]),
        .I1(\a9/k4a [9]),
        .O(k8b[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [0]),
        .Q(s1[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[100] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [100]),
        .Q(s1[100]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[101] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [101]),
        .Q(s1[101]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[102] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [102]),
        .Q(s1[102]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[103] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [103]),
        .Q(s1[103]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[104] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [104]),
        .Q(s1[104]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[105] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [105]),
        .Q(s1[105]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[106] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [106]),
        .Q(s1[106]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[107] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [107]),
        .Q(s1[107]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[108] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [108]),
        .Q(s1[108]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[109] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [109]),
        .Q(s1[109]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [10]),
        .Q(s1[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[110] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [110]),
        .Q(s1[110]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[111] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [111]),
        .Q(s1[111]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[112] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [112]),
        .Q(s1[112]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[113] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [113]),
        .Q(s1[113]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[114] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [114]),
        .Q(s1[114]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[115] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [115]),
        .Q(s1[115]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[116] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [116]),
        .Q(s1[116]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[117] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [117]),
        .Q(s1[117]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[118] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [118]),
        .Q(s1[118]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[119] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [119]),
        .Q(s1[119]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [11]),
        .Q(s1[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[120] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [120]),
        .Q(s1[120]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[121] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [121]),
        .Q(s1[121]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[122] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [122]),
        .Q(s1[122]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[123] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [123]),
        .Q(s1[123]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[124] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [124]),
        .Q(s1[124]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[125] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [125]),
        .Q(s1[125]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[126] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [126]),
        .Q(s1[126]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[127] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [127]),
        .Q(s1[127]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [12]),
        .Q(s1[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [13]),
        .Q(s1[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [14]),
        .Q(s1[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [15]),
        .Q(s1[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [16]),
        .Q(s1[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [17]),
        .Q(s1[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [18]),
        .Q(s1[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [19]),
        .Q(s1[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [1]),
        .Q(s1[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [20]),
        .Q(s1[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [21]),
        .Q(s1[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [22]),
        .Q(s1[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [23]),
        .Q(s1[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [24]),
        .Q(s1[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [25]),
        .Q(s1[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [26]),
        .Q(s1[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [27]),
        .Q(s1[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [28]),
        .Q(s1[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [29]),
        .Q(s1[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [2]),
        .Q(s1[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [30]),
        .Q(s1[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [31]),
        .Q(s1[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [32]),
        .Q(s1[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [33]),
        .Q(s1[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [34]),
        .Q(s1[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [35]),
        .Q(s1[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [36]),
        .Q(s1[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [37]),
        .Q(s1[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [38]),
        .Q(s1[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [39]),
        .Q(s1[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [3]),
        .Q(s1[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [40]),
        .Q(s1[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [41]),
        .Q(s1[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [42]),
        .Q(s1[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [43]),
        .Q(s1[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [44]),
        .Q(s1[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [45]),
        .Q(s1[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [46]),
        .Q(s1[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [47]),
        .Q(s1[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [48]),
        .Q(s1[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [49]),
        .Q(s1[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [4]),
        .Q(s1[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [50]),
        .Q(s1[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [51]),
        .Q(s1[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [52]),
        .Q(s1[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [53]),
        .Q(s1[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [54]),
        .Q(s1[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [55]),
        .Q(s1[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [56]),
        .Q(s1[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [57]),
        .Q(s1[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [58]),
        .Q(s1[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [59]),
        .Q(s1[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [5]),
        .Q(s1[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [60]),
        .Q(s1[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [61]),
        .Q(s1[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [62]),
        .Q(s1[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [63]),
        .Q(s1[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[64] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [64]),
        .Q(s1[64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[65] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [65]),
        .Q(s1[65]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[66] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [66]),
        .Q(s1[66]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[67] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [67]),
        .Q(s1[67]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[68] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [68]),
        .Q(s1[68]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[69] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [69]),
        .Q(s1[69]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [6]),
        .Q(s1[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[70] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [70]),
        .Q(s1[70]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[71] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [71]),
        .Q(s1[71]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[72] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [72]),
        .Q(s1[72]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[73] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [73]),
        .Q(s1[73]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[74] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [74]),
        .Q(s1[74]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[75] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [75]),
        .Q(s1[75]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[76] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [76]),
        .Q(s1[76]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[77] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [77]),
        .Q(s1[77]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[78] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [78]),
        .Q(s1[78]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[79] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [79]),
        .Q(s1[79]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [7]),
        .Q(s1[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[80] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [80]),
        .Q(s1[80]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[81] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [81]),
        .Q(s1[81]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[82] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [82]),
        .Q(s1[82]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[83] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [83]),
        .Q(s1[83]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[84] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [84]),
        .Q(s1[84]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[85] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [85]),
        .Q(s1[85]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[86] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [86]),
        .Q(s1[86]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[87] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [87]),
        .Q(s1[87]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[88] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [88]),
        .Q(s1[88]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[89] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [89]),
        .Q(s1[89]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [8]),
        .Q(s1[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[90] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [90]),
        .Q(s1[90]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[91] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [91]),
        .Q(s1[91]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[92] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [92]),
        .Q(s1[92]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[93] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [93]),
        .Q(s1[93]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[94] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [94]),
        .Q(s1[94]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[95] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [95]),
        .Q(s1[95]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[96] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [96]),
        .Q(s1[96]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[97] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [97]),
        .Q(s1[97]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[98] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [98]),
        .Q(s1[98]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[99] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [99]),
        .Q(s1[99]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r1/state_out_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r1/p_0_out [9]),
        .Q(s1[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r1/t0/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[127:120],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[119:112],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r1/t0/t0/s0/out_reg_n_0 ,\r1/t0/t0/s0/out_reg_n_1 ,\r1/t0/t0/s0/out_reg_n_2 ,\r1/t0/t0/s0/out_reg_n_3 ,\r1/t0/t0/s0/out_reg_n_4 ,\r1/t0/t0/s0/out_reg_n_5 ,\r1/t0/t0/s0/out_reg_n_6 ,\r1/t0/t0/s0/out_reg_n_7 ,\r1/t0/t0/p_0_in }),
        .DOBDO({\r1/t0/t0/s0/out_reg_n_16 ,\r1/t0/t0/s0/out_reg_n_17 ,\r1/t0/t0/s0/out_reg_n_18 ,\r1/t0/t0/s0/out_reg_n_19 ,\r1/t0/t0/s0/out_reg_n_20 ,\r1/t0/t0/s0/out_reg_n_21 ,\r1/t0/t0/s0/out_reg_n_22 ,\r1/t0/t0/s0/out_reg_n_23 ,\r1/t0/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r1/t0/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[127:120],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[119:112],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r1/t0/t0/s4/out_reg_n_0 ,\r1/t0/t0/s4/out_reg_n_1 ,\r1/t0/t0/s4/out_reg_n_2 ,\r1/t0/t0/s4/out_reg_n_3 ,\r1/t0/t0/s4/out_reg_n_4 ,\r1/t0/t0/s4/out_reg_n_5 ,\r1/t0/t0/s4/out_reg_n_6 ,\r1/t0/t0/s4/out_reg_n_7 ,\r1/t0/t0/p_1_in }),
        .DOBDO({\r1/t0/t0/s4/out_reg_n_16 ,\r1/t0/t0/s4/out_reg_n_17 ,\r1/t0/t0/s4/out_reg_n_18 ,\r1/t0/t0/s4/out_reg_n_19 ,\r1/t0/t0/s4/out_reg_n_20 ,\r1/t0/t0/s4/out_reg_n_21 ,\r1/t0/t0/s4/out_reg_n_22 ,\r1/t0/t0/s4/out_reg_n_23 ,\r1/t0/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r1/t0/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[111:104],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[103:96],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r1/t0/t2/s0/out_reg_n_0 ,\r1/t0/t2/s0/out_reg_n_1 ,\r1/t0/t2/s0/out_reg_n_2 ,\r1/t0/t2/s0/out_reg_n_3 ,\r1/t0/t2/s0/out_reg_n_4 ,\r1/t0/t2/s0/out_reg_n_5 ,\r1/t0/t2/s0/out_reg_n_6 ,\r1/t0/t2/s0/out_reg_n_7 ,\r1/t0/t2/p_0_in }),
        .DOBDO({\r1/t0/t2/s0/out_reg_n_16 ,\r1/t0/t2/s0/out_reg_n_17 ,\r1/t0/t2/s0/out_reg_n_18 ,\r1/t0/t2/s0/out_reg_n_19 ,\r1/t0/t2/s0/out_reg_n_20 ,\r1/t0/t2/s0/out_reg_n_21 ,\r1/t0/t2/s0/out_reg_n_22 ,\r1/t0/t2/s0/out_reg_n_23 ,\r1/t0/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r1/t0/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[111:104],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[103:96],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r1/t0/t2/s4/out_reg_n_0 ,\r1/t0/t2/s4/out_reg_n_1 ,\r1/t0/t2/s4/out_reg_n_2 ,\r1/t0/t2/s4/out_reg_n_3 ,\r1/t0/t2/s4/out_reg_n_4 ,\r1/t0/t2/s4/out_reg_n_5 ,\r1/t0/t2/s4/out_reg_n_6 ,\r1/t0/t2/s4/out_reg_n_7 ,\r1/t0/t2/p_1_in }),
        .DOBDO({\r1/t0/t2/s4/out_reg_n_16 ,\r1/t0/t2/s4/out_reg_n_17 ,\r1/t0/t2/s4/out_reg_n_18 ,\r1/t0/t2/s4/out_reg_n_19 ,\r1/t0/t2/s4/out_reg_n_20 ,\r1/t0/t2/s4/out_reg_n_21 ,\r1/t0/t2/s4/out_reg_n_22 ,\r1/t0/t2/s4/out_reg_n_23 ,\r1/t0/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r1/t1/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[95:88],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[87:80],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r1/t1/t0/s0/out_reg_n_0 ,\r1/t1/t0/s0/out_reg_n_1 ,\r1/t1/t0/s0/out_reg_n_2 ,\r1/t1/t0/s0/out_reg_n_3 ,\r1/t1/t0/s0/out_reg_n_4 ,\r1/t1/t0/s0/out_reg_n_5 ,\r1/t1/t0/s0/out_reg_n_6 ,\r1/t1/t0/s0/out_reg_n_7 ,\r1/t1/t0/p_0_in }),
        .DOBDO({\r1/t1/t0/s0/out_reg_n_16 ,\r1/t1/t0/s0/out_reg_n_17 ,\r1/t1/t0/s0/out_reg_n_18 ,\r1/t1/t0/s0/out_reg_n_19 ,\r1/t1/t0/s0/out_reg_n_20 ,\r1/t1/t0/s0/out_reg_n_21 ,\r1/t1/t0/s0/out_reg_n_22 ,\r1/t1/t0/s0/out_reg_n_23 ,\r1/t1/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r1/t1/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[95:88],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[87:80],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r1/t1/t0/s4/out_reg_n_0 ,\r1/t1/t0/s4/out_reg_n_1 ,\r1/t1/t0/s4/out_reg_n_2 ,\r1/t1/t0/s4/out_reg_n_3 ,\r1/t1/t0/s4/out_reg_n_4 ,\r1/t1/t0/s4/out_reg_n_5 ,\r1/t1/t0/s4/out_reg_n_6 ,\r1/t1/t0/s4/out_reg_n_7 ,\r1/t1/t0/p_1_in }),
        .DOBDO({\r1/t1/t0/s4/out_reg_n_16 ,\r1/t1/t0/s4/out_reg_n_17 ,\r1/t1/t0/s4/out_reg_n_18 ,\r1/t1/t0/s4/out_reg_n_19 ,\r1/t1/t0/s4/out_reg_n_20 ,\r1/t1/t0/s4/out_reg_n_21 ,\r1/t1/t0/s4/out_reg_n_22 ,\r1/t1/t0/s4/out_reg_n_23 ,\r1/t1/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r1/t1/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[79:72],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[71:64],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r1/t1/t2/s0/out_reg_n_0 ,\r1/t1/t2/s0/out_reg_n_1 ,\r1/t1/t2/s0/out_reg_n_2 ,\r1/t1/t2/s0/out_reg_n_3 ,\r1/t1/t2/s0/out_reg_n_4 ,\r1/t1/t2/s0/out_reg_n_5 ,\r1/t1/t2/s0/out_reg_n_6 ,\r1/t1/t2/s0/out_reg_n_7 ,\r1/t1/t2/p_0_in }),
        .DOBDO({\r1/t1/t2/s0/out_reg_n_16 ,\r1/t1/t2/s0/out_reg_n_17 ,\r1/t1/t2/s0/out_reg_n_18 ,\r1/t1/t2/s0/out_reg_n_19 ,\r1/t1/t2/s0/out_reg_n_20 ,\r1/t1/t2/s0/out_reg_n_21 ,\r1/t1/t2/s0/out_reg_n_22 ,\r1/t1/t2/s0/out_reg_n_23 ,\r1/t1/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r1/t1/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[79:72],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[71:64],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r1/t1/t2/s4/out_reg_n_0 ,\r1/t1/t2/s4/out_reg_n_1 ,\r1/t1/t2/s4/out_reg_n_2 ,\r1/t1/t2/s4/out_reg_n_3 ,\r1/t1/t2/s4/out_reg_n_4 ,\r1/t1/t2/s4/out_reg_n_5 ,\r1/t1/t2/s4/out_reg_n_6 ,\r1/t1/t2/s4/out_reg_n_7 ,\r1/t1/t2/p_1_in }),
        .DOBDO({\r1/t1/t2/s4/out_reg_n_16 ,\r1/t1/t2/s4/out_reg_n_17 ,\r1/t1/t2/s4/out_reg_n_18 ,\r1/t1/t2/s4/out_reg_n_19 ,\r1/t1/t2/s4/out_reg_n_20 ,\r1/t1/t2/s4/out_reg_n_21 ,\r1/t1/t2/s4/out_reg_n_22 ,\r1/t1/t2/s4/out_reg_n_23 ,\r1/t1/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r1/t2/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[63:56],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[55:48],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r1/t2/t0/s0/out_reg_n_0 ,\r1/t2/t0/s0/out_reg_n_1 ,\r1/t2/t0/s0/out_reg_n_2 ,\r1/t2/t0/s0/out_reg_n_3 ,\r1/t2/t0/s0/out_reg_n_4 ,\r1/t2/t0/s0/out_reg_n_5 ,\r1/t2/t0/s0/out_reg_n_6 ,\r1/t2/t0/s0/out_reg_n_7 ,\r1/t2/t0/p_0_in }),
        .DOBDO({\r1/t2/t0/s0/out_reg_n_16 ,\r1/t2/t0/s0/out_reg_n_17 ,\r1/t2/t0/s0/out_reg_n_18 ,\r1/t2/t0/s0/out_reg_n_19 ,\r1/t2/t0/s0/out_reg_n_20 ,\r1/t2/t0/s0/out_reg_n_21 ,\r1/t2/t0/s0/out_reg_n_22 ,\r1/t2/t0/s0/out_reg_n_23 ,\r1/t2/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r1/t2/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[63:56],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[55:48],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r1/t2/t0/s4/out_reg_n_0 ,\r1/t2/t0/s4/out_reg_n_1 ,\r1/t2/t0/s4/out_reg_n_2 ,\r1/t2/t0/s4/out_reg_n_3 ,\r1/t2/t0/s4/out_reg_n_4 ,\r1/t2/t0/s4/out_reg_n_5 ,\r1/t2/t0/s4/out_reg_n_6 ,\r1/t2/t0/s4/out_reg_n_7 ,\r1/t2/t0/p_1_in }),
        .DOBDO({\r1/t2/t0/s4/out_reg_n_16 ,\r1/t2/t0/s4/out_reg_n_17 ,\r1/t2/t0/s4/out_reg_n_18 ,\r1/t2/t0/s4/out_reg_n_19 ,\r1/t2/t0/s4/out_reg_n_20 ,\r1/t2/t0/s4/out_reg_n_21 ,\r1/t2/t0/s4/out_reg_n_22 ,\r1/t2/t0/s4/out_reg_n_23 ,\r1/t2/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r1/t2/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[47:40],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[39:32],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r1/t2/t2/s0/out_reg_n_0 ,\r1/t2/t2/s0/out_reg_n_1 ,\r1/t2/t2/s0/out_reg_n_2 ,\r1/t2/t2/s0/out_reg_n_3 ,\r1/t2/t2/s0/out_reg_n_4 ,\r1/t2/t2/s0/out_reg_n_5 ,\r1/t2/t2/s0/out_reg_n_6 ,\r1/t2/t2/s0/out_reg_n_7 ,\r1/t2/t2/p_0_in }),
        .DOBDO({\r1/t2/t2/s0/out_reg_n_16 ,\r1/t2/t2/s0/out_reg_n_17 ,\r1/t2/t2/s0/out_reg_n_18 ,\r1/t2/t2/s0/out_reg_n_19 ,\r1/t2/t2/s0/out_reg_n_20 ,\r1/t2/t2/s0/out_reg_n_21 ,\r1/t2/t2/s0/out_reg_n_22 ,\r1/t2/t2/s0/out_reg_n_23 ,\r1/t2/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r1/t2/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[47:40],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[39:32],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r1/t2/t2/s4/out_reg_n_0 ,\r1/t2/t2/s4/out_reg_n_1 ,\r1/t2/t2/s4/out_reg_n_2 ,\r1/t2/t2/s4/out_reg_n_3 ,\r1/t2/t2/s4/out_reg_n_4 ,\r1/t2/t2/s4/out_reg_n_5 ,\r1/t2/t2/s4/out_reg_n_6 ,\r1/t2/t2/s4/out_reg_n_7 ,\r1/t2/t2/p_1_in }),
        .DOBDO({\r1/t2/t2/s4/out_reg_n_16 ,\r1/t2/t2/s4/out_reg_n_17 ,\r1/t2/t2/s4/out_reg_n_18 ,\r1/t2/t2/s4/out_reg_n_19 ,\r1/t2/t2/s4/out_reg_n_20 ,\r1/t2/t2/s4/out_reg_n_21 ,\r1/t2/t2/s4/out_reg_n_22 ,\r1/t2/t2/s4/out_reg_n_23 ,\r1/t2/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r1/t3/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r1/t3/t0/s0/out_reg_n_0 ,\r1/t3/t0/s0/out_reg_n_1 ,\r1/t3/t0/s0/out_reg_n_2 ,\r1/t3/t0/s0/out_reg_n_3 ,\r1/t3/t0/s0/out_reg_n_4 ,\r1/t3/t0/s0/out_reg_n_5 ,\r1/t3/t0/s0/out_reg_n_6 ,\r1/t3/t0/s0/out_reg_n_7 ,\r1/t3/t0/p_0_in }),
        .DOBDO({\r1/t3/t0/s0/out_reg_n_16 ,\r1/t3/t0/s0/out_reg_n_17 ,\r1/t3/t0/s0/out_reg_n_18 ,\r1/t3/t0/s0/out_reg_n_19 ,\r1/t3/t0/s0/out_reg_n_20 ,\r1/t3/t0/s0/out_reg_n_21 ,\r1/t3/t0/s0/out_reg_n_22 ,\r1/t3/t0/s0/out_reg_n_23 ,\r1/t3/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r1/t3/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r1/t3/t0/s4/out_reg_n_0 ,\r1/t3/t0/s4/out_reg_n_1 ,\r1/t3/t0/s4/out_reg_n_2 ,\r1/t3/t0/s4/out_reg_n_3 ,\r1/t3/t0/s4/out_reg_n_4 ,\r1/t3/t0/s4/out_reg_n_5 ,\r1/t3/t0/s4/out_reg_n_6 ,\r1/t3/t0/s4/out_reg_n_7 ,\r1/t3/t0/p_1_in }),
        .DOBDO({\r1/t3/t0/s4/out_reg_n_16 ,\r1/t3/t0/s4/out_reg_n_17 ,\r1/t3/t0/s4/out_reg_n_18 ,\r1/t3/t0/s4/out_reg_n_19 ,\r1/t3/t0/s4/out_reg_n_20 ,\r1/t3/t0/s4/out_reg_n_21 ,\r1/t3/t0/s4/out_reg_n_22 ,\r1/t3/t0/s4/out_reg_n_23 ,\r1/t3/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r1/t3/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r1/t3/t2/s0/out_reg_n_0 ,\r1/t3/t2/s0/out_reg_n_1 ,\r1/t3/t2/s0/out_reg_n_2 ,\r1/t3/t2/s0/out_reg_n_3 ,\r1/t3/t2/s0/out_reg_n_4 ,\r1/t3/t2/s0/out_reg_n_5 ,\r1/t3/t2/s0/out_reg_n_6 ,\r1/t3/t2/s0/out_reg_n_7 ,\r1/t3/t2/p_0_in }),
        .DOBDO({\r1/t3/t2/s0/out_reg_n_16 ,\r1/t3/t2/s0/out_reg_n_17 ,\r1/t3/t2/s0/out_reg_n_18 ,\r1/t3/t2/s0/out_reg_n_19 ,\r1/t3/t2/s0/out_reg_n_20 ,\r1/t3/t2/s0/out_reg_n_21 ,\r1/t3/t2/s0/out_reg_n_22 ,\r1/t3/t2/s0/out_reg_n_23 ,\r1/t3/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r1/t3/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s0[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r1/t3/t2/s4/out_reg_n_0 ,\r1/t3/t2/s4/out_reg_n_1 ,\r1/t3/t2/s4/out_reg_n_2 ,\r1/t3/t2/s4/out_reg_n_3 ,\r1/t3/t2/s4/out_reg_n_4 ,\r1/t3/t2/s4/out_reg_n_5 ,\r1/t3/t2/s4/out_reg_n_6 ,\r1/t3/t2/s4/out_reg_n_7 ,\r1/t3/t2/p_1_in }),
        .DOBDO({\r1/t3/t2/s4/out_reg_n_16 ,\r1/t3/t2/s4/out_reg_n_17 ,\r1/t3/t2/s4/out_reg_n_18 ,\r1/t3/t2/s4/out_reg_n_19 ,\r1/t3/t2/s4/out_reg_n_20 ,\r1/t3/t2/s4/out_reg_n_21 ,\r1/t3/t2/s4/out_reg_n_22 ,\r1/t3/t2/s4/out_reg_n_23 ,\r1/t3/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [0]),
        .Q(s2[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[100] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [100]),
        .Q(s2[100]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[101] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [101]),
        .Q(s2[101]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[102] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [102]),
        .Q(s2[102]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[103] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [103]),
        .Q(s2[103]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[104] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [104]),
        .Q(s2[104]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[105] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [105]),
        .Q(s2[105]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[106] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [106]),
        .Q(s2[106]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[107] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [107]),
        .Q(s2[107]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[108] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [108]),
        .Q(s2[108]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[109] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [109]),
        .Q(s2[109]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [10]),
        .Q(s2[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[110] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [110]),
        .Q(s2[110]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[111] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [111]),
        .Q(s2[111]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[112] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [112]),
        .Q(s2[112]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[113] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [113]),
        .Q(s2[113]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[114] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [114]),
        .Q(s2[114]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[115] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [115]),
        .Q(s2[115]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[116] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [116]),
        .Q(s2[116]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[117] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [117]),
        .Q(s2[117]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[118] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [118]),
        .Q(s2[118]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[119] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [119]),
        .Q(s2[119]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [11]),
        .Q(s2[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[120] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [120]),
        .Q(s2[120]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[121] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [121]),
        .Q(s2[121]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[122] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [122]),
        .Q(s2[122]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[123] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [123]),
        .Q(s2[123]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[124] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [124]),
        .Q(s2[124]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[125] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [125]),
        .Q(s2[125]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[126] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [126]),
        .Q(s2[126]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[127] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [127]),
        .Q(s2[127]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [12]),
        .Q(s2[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [13]),
        .Q(s2[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [14]),
        .Q(s2[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [15]),
        .Q(s2[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [16]),
        .Q(s2[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [17]),
        .Q(s2[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [18]),
        .Q(s2[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [19]),
        .Q(s2[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [1]),
        .Q(s2[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [20]),
        .Q(s2[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [21]),
        .Q(s2[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [22]),
        .Q(s2[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [23]),
        .Q(s2[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [24]),
        .Q(s2[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [25]),
        .Q(s2[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [26]),
        .Q(s2[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [27]),
        .Q(s2[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [28]),
        .Q(s2[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [29]),
        .Q(s2[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [2]),
        .Q(s2[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [30]),
        .Q(s2[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [31]),
        .Q(s2[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [32]),
        .Q(s2[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [33]),
        .Q(s2[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [34]),
        .Q(s2[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [35]),
        .Q(s2[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [36]),
        .Q(s2[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [37]),
        .Q(s2[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [38]),
        .Q(s2[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [39]),
        .Q(s2[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [3]),
        .Q(s2[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [40]),
        .Q(s2[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [41]),
        .Q(s2[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [42]),
        .Q(s2[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [43]),
        .Q(s2[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [44]),
        .Q(s2[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [45]),
        .Q(s2[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [46]),
        .Q(s2[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [47]),
        .Q(s2[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [48]),
        .Q(s2[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [49]),
        .Q(s2[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [4]),
        .Q(s2[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [50]),
        .Q(s2[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [51]),
        .Q(s2[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [52]),
        .Q(s2[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [53]),
        .Q(s2[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [54]),
        .Q(s2[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [55]),
        .Q(s2[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [56]),
        .Q(s2[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [57]),
        .Q(s2[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [58]),
        .Q(s2[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [59]),
        .Q(s2[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [5]),
        .Q(s2[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [60]),
        .Q(s2[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [61]),
        .Q(s2[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [62]),
        .Q(s2[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [63]),
        .Q(s2[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[64] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [64]),
        .Q(s2[64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[65] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [65]),
        .Q(s2[65]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[66] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [66]),
        .Q(s2[66]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[67] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [67]),
        .Q(s2[67]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[68] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [68]),
        .Q(s2[68]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[69] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [69]),
        .Q(s2[69]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [6]),
        .Q(s2[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[70] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [70]),
        .Q(s2[70]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[71] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [71]),
        .Q(s2[71]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[72] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [72]),
        .Q(s2[72]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[73] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [73]),
        .Q(s2[73]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[74] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [74]),
        .Q(s2[74]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[75] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [75]),
        .Q(s2[75]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[76] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [76]),
        .Q(s2[76]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[77] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [77]),
        .Q(s2[77]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[78] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [78]),
        .Q(s2[78]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[79] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [79]),
        .Q(s2[79]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [7]),
        .Q(s2[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[80] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [80]),
        .Q(s2[80]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[81] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [81]),
        .Q(s2[81]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[82] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [82]),
        .Q(s2[82]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[83] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [83]),
        .Q(s2[83]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[84] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [84]),
        .Q(s2[84]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[85] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [85]),
        .Q(s2[85]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[86] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [86]),
        .Q(s2[86]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[87] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [87]),
        .Q(s2[87]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[88] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [88]),
        .Q(s2[88]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[89] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [89]),
        .Q(s2[89]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [8]),
        .Q(s2[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[90] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [90]),
        .Q(s2[90]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[91] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [91]),
        .Q(s2[91]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[92] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [92]),
        .Q(s2[92]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[93] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [93]),
        .Q(s2[93]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[94] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [94]),
        .Q(s2[94]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[95] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [95]),
        .Q(s2[95]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[96] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [96]),
        .Q(s2[96]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[97] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [97]),
        .Q(s2[97]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[98] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [98]),
        .Q(s2[98]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[99] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [99]),
        .Q(s2[99]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r2/state_out_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r2/p_0_out [9]),
        .Q(s2[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r2/t0/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[127:120],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[119:112],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r2/t0/t0/s0/out_reg_n_0 ,\r2/t0/t0/s0/out_reg_n_1 ,\r2/t0/t0/s0/out_reg_n_2 ,\r2/t0/t0/s0/out_reg_n_3 ,\r2/t0/t0/s0/out_reg_n_4 ,\r2/t0/t0/s0/out_reg_n_5 ,\r2/t0/t0/s0/out_reg_n_6 ,\r2/t0/t0/s0/out_reg_n_7 ,\r2/t0/t0/p_0_in }),
        .DOBDO({\r2/t0/t0/s0/out_reg_n_16 ,\r2/t0/t0/s0/out_reg_n_17 ,\r2/t0/t0/s0/out_reg_n_18 ,\r2/t0/t0/s0/out_reg_n_19 ,\r2/t0/t0/s0/out_reg_n_20 ,\r2/t0/t0/s0/out_reg_n_21 ,\r2/t0/t0/s0/out_reg_n_22 ,\r2/t0/t0/s0/out_reg_n_23 ,\r2/t0/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r2/t0/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[127:120],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[119:112],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r2/t0/t0/s4/out_reg_n_0 ,\r2/t0/t0/s4/out_reg_n_1 ,\r2/t0/t0/s4/out_reg_n_2 ,\r2/t0/t0/s4/out_reg_n_3 ,\r2/t0/t0/s4/out_reg_n_4 ,\r2/t0/t0/s4/out_reg_n_5 ,\r2/t0/t0/s4/out_reg_n_6 ,\r2/t0/t0/s4/out_reg_n_7 ,\r2/t0/t0/p_1_in }),
        .DOBDO({\r2/t0/t0/s4/out_reg_n_16 ,\r2/t0/t0/s4/out_reg_n_17 ,\r2/t0/t0/s4/out_reg_n_18 ,\r2/t0/t0/s4/out_reg_n_19 ,\r2/t0/t0/s4/out_reg_n_20 ,\r2/t0/t0/s4/out_reg_n_21 ,\r2/t0/t0/s4/out_reg_n_22 ,\r2/t0/t0/s4/out_reg_n_23 ,\r2/t0/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r2/t0/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[111:104],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[103:96],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r2/t0/t2/s0/out_reg_n_0 ,\r2/t0/t2/s0/out_reg_n_1 ,\r2/t0/t2/s0/out_reg_n_2 ,\r2/t0/t2/s0/out_reg_n_3 ,\r2/t0/t2/s0/out_reg_n_4 ,\r2/t0/t2/s0/out_reg_n_5 ,\r2/t0/t2/s0/out_reg_n_6 ,\r2/t0/t2/s0/out_reg_n_7 ,\r2/t0/t2/p_0_in }),
        .DOBDO({\r2/t0/t2/s0/out_reg_n_16 ,\r2/t0/t2/s0/out_reg_n_17 ,\r2/t0/t2/s0/out_reg_n_18 ,\r2/t0/t2/s0/out_reg_n_19 ,\r2/t0/t2/s0/out_reg_n_20 ,\r2/t0/t2/s0/out_reg_n_21 ,\r2/t0/t2/s0/out_reg_n_22 ,\r2/t0/t2/s0/out_reg_n_23 ,\r2/t0/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r2/t0/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[111:104],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[103:96],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r2/t0/t2/s4/out_reg_n_0 ,\r2/t0/t2/s4/out_reg_n_1 ,\r2/t0/t2/s4/out_reg_n_2 ,\r2/t0/t2/s4/out_reg_n_3 ,\r2/t0/t2/s4/out_reg_n_4 ,\r2/t0/t2/s4/out_reg_n_5 ,\r2/t0/t2/s4/out_reg_n_6 ,\r2/t0/t2/s4/out_reg_n_7 ,\r2/t0/t2/p_1_in }),
        .DOBDO({\r2/t0/t2/s4/out_reg_n_16 ,\r2/t0/t2/s4/out_reg_n_17 ,\r2/t0/t2/s4/out_reg_n_18 ,\r2/t0/t2/s4/out_reg_n_19 ,\r2/t0/t2/s4/out_reg_n_20 ,\r2/t0/t2/s4/out_reg_n_21 ,\r2/t0/t2/s4/out_reg_n_22 ,\r2/t0/t2/s4/out_reg_n_23 ,\r2/t0/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r2/t1/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[95:88],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[87:80],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r2/t1/t0/s0/out_reg_n_0 ,\r2/t1/t0/s0/out_reg_n_1 ,\r2/t1/t0/s0/out_reg_n_2 ,\r2/t1/t0/s0/out_reg_n_3 ,\r2/t1/t0/s0/out_reg_n_4 ,\r2/t1/t0/s0/out_reg_n_5 ,\r2/t1/t0/s0/out_reg_n_6 ,\r2/t1/t0/s0/out_reg_n_7 ,\r2/t1/t0/p_0_in }),
        .DOBDO({\r2/t1/t0/s0/out_reg_n_16 ,\r2/t1/t0/s0/out_reg_n_17 ,\r2/t1/t0/s0/out_reg_n_18 ,\r2/t1/t0/s0/out_reg_n_19 ,\r2/t1/t0/s0/out_reg_n_20 ,\r2/t1/t0/s0/out_reg_n_21 ,\r2/t1/t0/s0/out_reg_n_22 ,\r2/t1/t0/s0/out_reg_n_23 ,\r2/t1/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r2/t1/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[95:88],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[87:80],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r2/t1/t0/s4/out_reg_n_0 ,\r2/t1/t0/s4/out_reg_n_1 ,\r2/t1/t0/s4/out_reg_n_2 ,\r2/t1/t0/s4/out_reg_n_3 ,\r2/t1/t0/s4/out_reg_n_4 ,\r2/t1/t0/s4/out_reg_n_5 ,\r2/t1/t0/s4/out_reg_n_6 ,\r2/t1/t0/s4/out_reg_n_7 ,\r2/t1/t0/p_1_in }),
        .DOBDO({\r2/t1/t0/s4/out_reg_n_16 ,\r2/t1/t0/s4/out_reg_n_17 ,\r2/t1/t0/s4/out_reg_n_18 ,\r2/t1/t0/s4/out_reg_n_19 ,\r2/t1/t0/s4/out_reg_n_20 ,\r2/t1/t0/s4/out_reg_n_21 ,\r2/t1/t0/s4/out_reg_n_22 ,\r2/t1/t0/s4/out_reg_n_23 ,\r2/t1/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r2/t1/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[79:72],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[71:64],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r2/t1/t2/s0/out_reg_n_0 ,\r2/t1/t2/s0/out_reg_n_1 ,\r2/t1/t2/s0/out_reg_n_2 ,\r2/t1/t2/s0/out_reg_n_3 ,\r2/t1/t2/s0/out_reg_n_4 ,\r2/t1/t2/s0/out_reg_n_5 ,\r2/t1/t2/s0/out_reg_n_6 ,\r2/t1/t2/s0/out_reg_n_7 ,\r2/t1/t2/p_0_in }),
        .DOBDO({\r2/t1/t2/s0/out_reg_n_16 ,\r2/t1/t2/s0/out_reg_n_17 ,\r2/t1/t2/s0/out_reg_n_18 ,\r2/t1/t2/s0/out_reg_n_19 ,\r2/t1/t2/s0/out_reg_n_20 ,\r2/t1/t2/s0/out_reg_n_21 ,\r2/t1/t2/s0/out_reg_n_22 ,\r2/t1/t2/s0/out_reg_n_23 ,\r2/t1/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r2/t1/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[79:72],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[71:64],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r2/t1/t2/s4/out_reg_n_0 ,\r2/t1/t2/s4/out_reg_n_1 ,\r2/t1/t2/s4/out_reg_n_2 ,\r2/t1/t2/s4/out_reg_n_3 ,\r2/t1/t2/s4/out_reg_n_4 ,\r2/t1/t2/s4/out_reg_n_5 ,\r2/t1/t2/s4/out_reg_n_6 ,\r2/t1/t2/s4/out_reg_n_7 ,\r2/t1/t2/p_1_in }),
        .DOBDO({\r2/t1/t2/s4/out_reg_n_16 ,\r2/t1/t2/s4/out_reg_n_17 ,\r2/t1/t2/s4/out_reg_n_18 ,\r2/t1/t2/s4/out_reg_n_19 ,\r2/t1/t2/s4/out_reg_n_20 ,\r2/t1/t2/s4/out_reg_n_21 ,\r2/t1/t2/s4/out_reg_n_22 ,\r2/t1/t2/s4/out_reg_n_23 ,\r2/t1/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r2/t2/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[63:56],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[55:48],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r2/t2/t0/s0/out_reg_n_0 ,\r2/t2/t0/s0/out_reg_n_1 ,\r2/t2/t0/s0/out_reg_n_2 ,\r2/t2/t0/s0/out_reg_n_3 ,\r2/t2/t0/s0/out_reg_n_4 ,\r2/t2/t0/s0/out_reg_n_5 ,\r2/t2/t0/s0/out_reg_n_6 ,\r2/t2/t0/s0/out_reg_n_7 ,\r2/t2/t0/p_0_in }),
        .DOBDO({\r2/t2/t0/s0/out_reg_n_16 ,\r2/t2/t0/s0/out_reg_n_17 ,\r2/t2/t0/s0/out_reg_n_18 ,\r2/t2/t0/s0/out_reg_n_19 ,\r2/t2/t0/s0/out_reg_n_20 ,\r2/t2/t0/s0/out_reg_n_21 ,\r2/t2/t0/s0/out_reg_n_22 ,\r2/t2/t0/s0/out_reg_n_23 ,\r2/t2/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r2/t2/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[63:56],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[55:48],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r2/t2/t0/s4/out_reg_n_0 ,\r2/t2/t0/s4/out_reg_n_1 ,\r2/t2/t0/s4/out_reg_n_2 ,\r2/t2/t0/s4/out_reg_n_3 ,\r2/t2/t0/s4/out_reg_n_4 ,\r2/t2/t0/s4/out_reg_n_5 ,\r2/t2/t0/s4/out_reg_n_6 ,\r2/t2/t0/s4/out_reg_n_7 ,\r2/t2/t0/p_1_in }),
        .DOBDO({\r2/t2/t0/s4/out_reg_n_16 ,\r2/t2/t0/s4/out_reg_n_17 ,\r2/t2/t0/s4/out_reg_n_18 ,\r2/t2/t0/s4/out_reg_n_19 ,\r2/t2/t0/s4/out_reg_n_20 ,\r2/t2/t0/s4/out_reg_n_21 ,\r2/t2/t0/s4/out_reg_n_22 ,\r2/t2/t0/s4/out_reg_n_23 ,\r2/t2/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r2/t2/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[47:40],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[39:32],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r2/t2/t2/s0/out_reg_n_0 ,\r2/t2/t2/s0/out_reg_n_1 ,\r2/t2/t2/s0/out_reg_n_2 ,\r2/t2/t2/s0/out_reg_n_3 ,\r2/t2/t2/s0/out_reg_n_4 ,\r2/t2/t2/s0/out_reg_n_5 ,\r2/t2/t2/s0/out_reg_n_6 ,\r2/t2/t2/s0/out_reg_n_7 ,\r2/t2/t2/p_0_in }),
        .DOBDO({\r2/t2/t2/s0/out_reg_n_16 ,\r2/t2/t2/s0/out_reg_n_17 ,\r2/t2/t2/s0/out_reg_n_18 ,\r2/t2/t2/s0/out_reg_n_19 ,\r2/t2/t2/s0/out_reg_n_20 ,\r2/t2/t2/s0/out_reg_n_21 ,\r2/t2/t2/s0/out_reg_n_22 ,\r2/t2/t2/s0/out_reg_n_23 ,\r2/t2/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r2/t2/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[47:40],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[39:32],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r2/t2/t2/s4/out_reg_n_0 ,\r2/t2/t2/s4/out_reg_n_1 ,\r2/t2/t2/s4/out_reg_n_2 ,\r2/t2/t2/s4/out_reg_n_3 ,\r2/t2/t2/s4/out_reg_n_4 ,\r2/t2/t2/s4/out_reg_n_5 ,\r2/t2/t2/s4/out_reg_n_6 ,\r2/t2/t2/s4/out_reg_n_7 ,\r2/t2/t2/p_1_in }),
        .DOBDO({\r2/t2/t2/s4/out_reg_n_16 ,\r2/t2/t2/s4/out_reg_n_17 ,\r2/t2/t2/s4/out_reg_n_18 ,\r2/t2/t2/s4/out_reg_n_19 ,\r2/t2/t2/s4/out_reg_n_20 ,\r2/t2/t2/s4/out_reg_n_21 ,\r2/t2/t2/s4/out_reg_n_22 ,\r2/t2/t2/s4/out_reg_n_23 ,\r2/t2/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r2/t3/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r2/t3/t0/s0/out_reg_n_0 ,\r2/t3/t0/s0/out_reg_n_1 ,\r2/t3/t0/s0/out_reg_n_2 ,\r2/t3/t0/s0/out_reg_n_3 ,\r2/t3/t0/s0/out_reg_n_4 ,\r2/t3/t0/s0/out_reg_n_5 ,\r2/t3/t0/s0/out_reg_n_6 ,\r2/t3/t0/s0/out_reg_n_7 ,\r2/t3/t0/p_0_in }),
        .DOBDO({\r2/t3/t0/s0/out_reg_n_16 ,\r2/t3/t0/s0/out_reg_n_17 ,\r2/t3/t0/s0/out_reg_n_18 ,\r2/t3/t0/s0/out_reg_n_19 ,\r2/t3/t0/s0/out_reg_n_20 ,\r2/t3/t0/s0/out_reg_n_21 ,\r2/t3/t0/s0/out_reg_n_22 ,\r2/t3/t0/s0/out_reg_n_23 ,\r2/t3/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r2/t3/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r2/t3/t0/s4/out_reg_n_0 ,\r2/t3/t0/s4/out_reg_n_1 ,\r2/t3/t0/s4/out_reg_n_2 ,\r2/t3/t0/s4/out_reg_n_3 ,\r2/t3/t0/s4/out_reg_n_4 ,\r2/t3/t0/s4/out_reg_n_5 ,\r2/t3/t0/s4/out_reg_n_6 ,\r2/t3/t0/s4/out_reg_n_7 ,\r2/t3/t0/p_1_in }),
        .DOBDO({\r2/t3/t0/s4/out_reg_n_16 ,\r2/t3/t0/s4/out_reg_n_17 ,\r2/t3/t0/s4/out_reg_n_18 ,\r2/t3/t0/s4/out_reg_n_19 ,\r2/t3/t0/s4/out_reg_n_20 ,\r2/t3/t0/s4/out_reg_n_21 ,\r2/t3/t0/s4/out_reg_n_22 ,\r2/t3/t0/s4/out_reg_n_23 ,\r2/t3/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r2/t3/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r2/t3/t2/s0/out_reg_n_0 ,\r2/t3/t2/s0/out_reg_n_1 ,\r2/t3/t2/s0/out_reg_n_2 ,\r2/t3/t2/s0/out_reg_n_3 ,\r2/t3/t2/s0/out_reg_n_4 ,\r2/t3/t2/s0/out_reg_n_5 ,\r2/t3/t2/s0/out_reg_n_6 ,\r2/t3/t2/s0/out_reg_n_7 ,\r2/t3/t2/p_0_in }),
        .DOBDO({\r2/t3/t2/s0/out_reg_n_16 ,\r2/t3/t2/s0/out_reg_n_17 ,\r2/t3/t2/s0/out_reg_n_18 ,\r2/t3/t2/s0/out_reg_n_19 ,\r2/t3/t2/s0/out_reg_n_20 ,\r2/t3/t2/s0/out_reg_n_21 ,\r2/t3/t2/s0/out_reg_n_22 ,\r2/t3/t2/s0/out_reg_n_23 ,\r2/t3/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r2/t3/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s1[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r2/t3/t2/s4/out_reg_n_0 ,\r2/t3/t2/s4/out_reg_n_1 ,\r2/t3/t2/s4/out_reg_n_2 ,\r2/t3/t2/s4/out_reg_n_3 ,\r2/t3/t2/s4/out_reg_n_4 ,\r2/t3/t2/s4/out_reg_n_5 ,\r2/t3/t2/s4/out_reg_n_6 ,\r2/t3/t2/s4/out_reg_n_7 ,\r2/t3/t2/p_1_in }),
        .DOBDO({\r2/t3/t2/s4/out_reg_n_16 ,\r2/t3/t2/s4/out_reg_n_17 ,\r2/t3/t2/s4/out_reg_n_18 ,\r2/t3/t2/s4/out_reg_n_19 ,\r2/t3/t2/s4/out_reg_n_20 ,\r2/t3/t2/s4/out_reg_n_21 ,\r2/t3/t2/s4/out_reg_n_22 ,\r2/t3/t2/s4/out_reg_n_23 ,\r2/t3/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [0]),
        .Q(s3[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[100] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [100]),
        .Q(s3[100]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[101] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [101]),
        .Q(s3[101]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[102] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [102]),
        .Q(s3[102]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[103] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [103]),
        .Q(s3[103]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[104] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [104]),
        .Q(s3[104]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[105] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [105]),
        .Q(s3[105]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[106] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [106]),
        .Q(s3[106]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[107] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [107]),
        .Q(s3[107]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[108] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [108]),
        .Q(s3[108]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[109] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [109]),
        .Q(s3[109]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [10]),
        .Q(s3[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[110] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [110]),
        .Q(s3[110]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[111] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [111]),
        .Q(s3[111]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[112] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [112]),
        .Q(s3[112]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[113] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [113]),
        .Q(s3[113]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[114] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [114]),
        .Q(s3[114]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[115] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [115]),
        .Q(s3[115]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[116] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [116]),
        .Q(s3[116]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[117] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [117]),
        .Q(s3[117]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[118] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [118]),
        .Q(s3[118]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[119] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [119]),
        .Q(s3[119]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [11]),
        .Q(s3[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[120] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [120]),
        .Q(s3[120]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[121] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [121]),
        .Q(s3[121]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[122] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [122]),
        .Q(s3[122]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[123] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [123]),
        .Q(s3[123]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[124] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [124]),
        .Q(s3[124]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[125] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [125]),
        .Q(s3[125]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[126] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [126]),
        .Q(s3[126]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[127] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [127]),
        .Q(s3[127]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [12]),
        .Q(s3[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [13]),
        .Q(s3[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [14]),
        .Q(s3[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [15]),
        .Q(s3[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [16]),
        .Q(s3[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [17]),
        .Q(s3[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [18]),
        .Q(s3[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [19]),
        .Q(s3[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [1]),
        .Q(s3[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [20]),
        .Q(s3[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [21]),
        .Q(s3[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [22]),
        .Q(s3[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [23]),
        .Q(s3[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [24]),
        .Q(s3[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [25]),
        .Q(s3[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [26]),
        .Q(s3[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [27]),
        .Q(s3[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [28]),
        .Q(s3[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [29]),
        .Q(s3[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [2]),
        .Q(s3[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [30]),
        .Q(s3[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [31]),
        .Q(s3[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [32]),
        .Q(s3[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [33]),
        .Q(s3[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [34]),
        .Q(s3[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [35]),
        .Q(s3[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [36]),
        .Q(s3[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [37]),
        .Q(s3[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [38]),
        .Q(s3[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [39]),
        .Q(s3[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [3]),
        .Q(s3[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [40]),
        .Q(s3[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [41]),
        .Q(s3[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [42]),
        .Q(s3[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [43]),
        .Q(s3[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [44]),
        .Q(s3[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [45]),
        .Q(s3[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [46]),
        .Q(s3[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [47]),
        .Q(s3[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [48]),
        .Q(s3[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [49]),
        .Q(s3[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [4]),
        .Q(s3[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [50]),
        .Q(s3[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [51]),
        .Q(s3[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [52]),
        .Q(s3[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [53]),
        .Q(s3[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [54]),
        .Q(s3[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [55]),
        .Q(s3[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [56]),
        .Q(s3[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [57]),
        .Q(s3[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [58]),
        .Q(s3[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [59]),
        .Q(s3[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [5]),
        .Q(s3[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [60]),
        .Q(s3[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [61]),
        .Q(s3[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [62]),
        .Q(s3[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [63]),
        .Q(s3[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[64] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [64]),
        .Q(s3[64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[65] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [65]),
        .Q(s3[65]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[66] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [66]),
        .Q(s3[66]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[67] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [67]),
        .Q(s3[67]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[68] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [68]),
        .Q(s3[68]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[69] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [69]),
        .Q(s3[69]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [6]),
        .Q(s3[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[70] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [70]),
        .Q(s3[70]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[71] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [71]),
        .Q(s3[71]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[72] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [72]),
        .Q(s3[72]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[73] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [73]),
        .Q(s3[73]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[74] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [74]),
        .Q(s3[74]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[75] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [75]),
        .Q(s3[75]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[76] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [76]),
        .Q(s3[76]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[77] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [77]),
        .Q(s3[77]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[78] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [78]),
        .Q(s3[78]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[79] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [79]),
        .Q(s3[79]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [7]),
        .Q(s3[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[80] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [80]),
        .Q(s3[80]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[81] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [81]),
        .Q(s3[81]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[82] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [82]),
        .Q(s3[82]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[83] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [83]),
        .Q(s3[83]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[84] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [84]),
        .Q(s3[84]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[85] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [85]),
        .Q(s3[85]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[86] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [86]),
        .Q(s3[86]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[87] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [87]),
        .Q(s3[87]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[88] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [88]),
        .Q(s3[88]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[89] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [89]),
        .Q(s3[89]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [8]),
        .Q(s3[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[90] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [90]),
        .Q(s3[90]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[91] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [91]),
        .Q(s3[91]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[92] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [92]),
        .Q(s3[92]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[93] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [93]),
        .Q(s3[93]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[94] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [94]),
        .Q(s3[94]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[95] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [95]),
        .Q(s3[95]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[96] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [96]),
        .Q(s3[96]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[97] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [97]),
        .Q(s3[97]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[98] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [98]),
        .Q(s3[98]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[99] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [99]),
        .Q(s3[99]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r3/state_out_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r3/p_0_out [9]),
        .Q(s3[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r3/t0/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[127:120],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[119:112],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r3/t0/t0/s0/out_reg_n_0 ,\r3/t0/t0/s0/out_reg_n_1 ,\r3/t0/t0/s0/out_reg_n_2 ,\r3/t0/t0/s0/out_reg_n_3 ,\r3/t0/t0/s0/out_reg_n_4 ,\r3/t0/t0/s0/out_reg_n_5 ,\r3/t0/t0/s0/out_reg_n_6 ,\r3/t0/t0/s0/out_reg_n_7 ,\r3/t0/t0/p_0_in }),
        .DOBDO({\r3/t0/t0/s0/out_reg_n_16 ,\r3/t0/t0/s0/out_reg_n_17 ,\r3/t0/t0/s0/out_reg_n_18 ,\r3/t0/t0/s0/out_reg_n_19 ,\r3/t0/t0/s0/out_reg_n_20 ,\r3/t0/t0/s0/out_reg_n_21 ,\r3/t0/t0/s0/out_reg_n_22 ,\r3/t0/t0/s0/out_reg_n_23 ,\r3/t0/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r3/t0/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[127:120],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[119:112],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r3/t0/t0/s4/out_reg_n_0 ,\r3/t0/t0/s4/out_reg_n_1 ,\r3/t0/t0/s4/out_reg_n_2 ,\r3/t0/t0/s4/out_reg_n_3 ,\r3/t0/t0/s4/out_reg_n_4 ,\r3/t0/t0/s4/out_reg_n_5 ,\r3/t0/t0/s4/out_reg_n_6 ,\r3/t0/t0/s4/out_reg_n_7 ,\r3/t0/t0/p_1_in }),
        .DOBDO({\r3/t0/t0/s4/out_reg_n_16 ,\r3/t0/t0/s4/out_reg_n_17 ,\r3/t0/t0/s4/out_reg_n_18 ,\r3/t0/t0/s4/out_reg_n_19 ,\r3/t0/t0/s4/out_reg_n_20 ,\r3/t0/t0/s4/out_reg_n_21 ,\r3/t0/t0/s4/out_reg_n_22 ,\r3/t0/t0/s4/out_reg_n_23 ,\r3/t0/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r3/t0/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[111:104],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[103:96],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r3/t0/t2/s0/out_reg_n_0 ,\r3/t0/t2/s0/out_reg_n_1 ,\r3/t0/t2/s0/out_reg_n_2 ,\r3/t0/t2/s0/out_reg_n_3 ,\r3/t0/t2/s0/out_reg_n_4 ,\r3/t0/t2/s0/out_reg_n_5 ,\r3/t0/t2/s0/out_reg_n_6 ,\r3/t0/t2/s0/out_reg_n_7 ,\r3/t0/t2/p_0_in }),
        .DOBDO({\r3/t0/t2/s0/out_reg_n_16 ,\r3/t0/t2/s0/out_reg_n_17 ,\r3/t0/t2/s0/out_reg_n_18 ,\r3/t0/t2/s0/out_reg_n_19 ,\r3/t0/t2/s0/out_reg_n_20 ,\r3/t0/t2/s0/out_reg_n_21 ,\r3/t0/t2/s0/out_reg_n_22 ,\r3/t0/t2/s0/out_reg_n_23 ,\r3/t0/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r3/t0/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[111:104],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[103:96],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r3/t0/t2/s4/out_reg_n_0 ,\r3/t0/t2/s4/out_reg_n_1 ,\r3/t0/t2/s4/out_reg_n_2 ,\r3/t0/t2/s4/out_reg_n_3 ,\r3/t0/t2/s4/out_reg_n_4 ,\r3/t0/t2/s4/out_reg_n_5 ,\r3/t0/t2/s4/out_reg_n_6 ,\r3/t0/t2/s4/out_reg_n_7 ,\r3/t0/t2/p_1_in }),
        .DOBDO({\r3/t0/t2/s4/out_reg_n_16 ,\r3/t0/t2/s4/out_reg_n_17 ,\r3/t0/t2/s4/out_reg_n_18 ,\r3/t0/t2/s4/out_reg_n_19 ,\r3/t0/t2/s4/out_reg_n_20 ,\r3/t0/t2/s4/out_reg_n_21 ,\r3/t0/t2/s4/out_reg_n_22 ,\r3/t0/t2/s4/out_reg_n_23 ,\r3/t0/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r3/t1/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[95:88],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[87:80],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r3/t1/t0/s0/out_reg_n_0 ,\r3/t1/t0/s0/out_reg_n_1 ,\r3/t1/t0/s0/out_reg_n_2 ,\r3/t1/t0/s0/out_reg_n_3 ,\r3/t1/t0/s0/out_reg_n_4 ,\r3/t1/t0/s0/out_reg_n_5 ,\r3/t1/t0/s0/out_reg_n_6 ,\r3/t1/t0/s0/out_reg_n_7 ,\r3/t1/t0/p_0_in }),
        .DOBDO({\r3/t1/t0/s0/out_reg_n_16 ,\r3/t1/t0/s0/out_reg_n_17 ,\r3/t1/t0/s0/out_reg_n_18 ,\r3/t1/t0/s0/out_reg_n_19 ,\r3/t1/t0/s0/out_reg_n_20 ,\r3/t1/t0/s0/out_reg_n_21 ,\r3/t1/t0/s0/out_reg_n_22 ,\r3/t1/t0/s0/out_reg_n_23 ,\r3/t1/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r3/t1/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[95:88],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[87:80],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r3/t1/t0/s4/out_reg_n_0 ,\r3/t1/t0/s4/out_reg_n_1 ,\r3/t1/t0/s4/out_reg_n_2 ,\r3/t1/t0/s4/out_reg_n_3 ,\r3/t1/t0/s4/out_reg_n_4 ,\r3/t1/t0/s4/out_reg_n_5 ,\r3/t1/t0/s4/out_reg_n_6 ,\r3/t1/t0/s4/out_reg_n_7 ,\r3/t1/t0/p_1_in }),
        .DOBDO({\r3/t1/t0/s4/out_reg_n_16 ,\r3/t1/t0/s4/out_reg_n_17 ,\r3/t1/t0/s4/out_reg_n_18 ,\r3/t1/t0/s4/out_reg_n_19 ,\r3/t1/t0/s4/out_reg_n_20 ,\r3/t1/t0/s4/out_reg_n_21 ,\r3/t1/t0/s4/out_reg_n_22 ,\r3/t1/t0/s4/out_reg_n_23 ,\r3/t1/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r3/t1/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[79:72],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[71:64],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r3/t1/t2/s0/out_reg_n_0 ,\r3/t1/t2/s0/out_reg_n_1 ,\r3/t1/t2/s0/out_reg_n_2 ,\r3/t1/t2/s0/out_reg_n_3 ,\r3/t1/t2/s0/out_reg_n_4 ,\r3/t1/t2/s0/out_reg_n_5 ,\r3/t1/t2/s0/out_reg_n_6 ,\r3/t1/t2/s0/out_reg_n_7 ,\r3/t1/t2/p_0_in }),
        .DOBDO({\r3/t1/t2/s0/out_reg_n_16 ,\r3/t1/t2/s0/out_reg_n_17 ,\r3/t1/t2/s0/out_reg_n_18 ,\r3/t1/t2/s0/out_reg_n_19 ,\r3/t1/t2/s0/out_reg_n_20 ,\r3/t1/t2/s0/out_reg_n_21 ,\r3/t1/t2/s0/out_reg_n_22 ,\r3/t1/t2/s0/out_reg_n_23 ,\r3/t1/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r3/t1/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[79:72],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[71:64],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r3/t1/t2/s4/out_reg_n_0 ,\r3/t1/t2/s4/out_reg_n_1 ,\r3/t1/t2/s4/out_reg_n_2 ,\r3/t1/t2/s4/out_reg_n_3 ,\r3/t1/t2/s4/out_reg_n_4 ,\r3/t1/t2/s4/out_reg_n_5 ,\r3/t1/t2/s4/out_reg_n_6 ,\r3/t1/t2/s4/out_reg_n_7 ,\r3/t1/t2/p_1_in }),
        .DOBDO({\r3/t1/t2/s4/out_reg_n_16 ,\r3/t1/t2/s4/out_reg_n_17 ,\r3/t1/t2/s4/out_reg_n_18 ,\r3/t1/t2/s4/out_reg_n_19 ,\r3/t1/t2/s4/out_reg_n_20 ,\r3/t1/t2/s4/out_reg_n_21 ,\r3/t1/t2/s4/out_reg_n_22 ,\r3/t1/t2/s4/out_reg_n_23 ,\r3/t1/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r3/t2/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[63:56],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[55:48],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r3/t2/t0/s0/out_reg_n_0 ,\r3/t2/t0/s0/out_reg_n_1 ,\r3/t2/t0/s0/out_reg_n_2 ,\r3/t2/t0/s0/out_reg_n_3 ,\r3/t2/t0/s0/out_reg_n_4 ,\r3/t2/t0/s0/out_reg_n_5 ,\r3/t2/t0/s0/out_reg_n_6 ,\r3/t2/t0/s0/out_reg_n_7 ,\r3/t2/t0/p_0_in }),
        .DOBDO({\r3/t2/t0/s0/out_reg_n_16 ,\r3/t2/t0/s0/out_reg_n_17 ,\r3/t2/t0/s0/out_reg_n_18 ,\r3/t2/t0/s0/out_reg_n_19 ,\r3/t2/t0/s0/out_reg_n_20 ,\r3/t2/t0/s0/out_reg_n_21 ,\r3/t2/t0/s0/out_reg_n_22 ,\r3/t2/t0/s0/out_reg_n_23 ,\r3/t2/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r3/t2/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[63:56],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[55:48],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r3/t2/t0/s4/out_reg_n_0 ,\r3/t2/t0/s4/out_reg_n_1 ,\r3/t2/t0/s4/out_reg_n_2 ,\r3/t2/t0/s4/out_reg_n_3 ,\r3/t2/t0/s4/out_reg_n_4 ,\r3/t2/t0/s4/out_reg_n_5 ,\r3/t2/t0/s4/out_reg_n_6 ,\r3/t2/t0/s4/out_reg_n_7 ,\r3/t2/t0/p_1_in }),
        .DOBDO({\r3/t2/t0/s4/out_reg_n_16 ,\r3/t2/t0/s4/out_reg_n_17 ,\r3/t2/t0/s4/out_reg_n_18 ,\r3/t2/t0/s4/out_reg_n_19 ,\r3/t2/t0/s4/out_reg_n_20 ,\r3/t2/t0/s4/out_reg_n_21 ,\r3/t2/t0/s4/out_reg_n_22 ,\r3/t2/t0/s4/out_reg_n_23 ,\r3/t2/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r3/t2/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[47:40],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[39:32],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r3/t2/t2/s0/out_reg_n_0 ,\r3/t2/t2/s0/out_reg_n_1 ,\r3/t2/t2/s0/out_reg_n_2 ,\r3/t2/t2/s0/out_reg_n_3 ,\r3/t2/t2/s0/out_reg_n_4 ,\r3/t2/t2/s0/out_reg_n_5 ,\r3/t2/t2/s0/out_reg_n_6 ,\r3/t2/t2/s0/out_reg_n_7 ,\r3/t2/t2/p_0_in }),
        .DOBDO({\r3/t2/t2/s0/out_reg_n_16 ,\r3/t2/t2/s0/out_reg_n_17 ,\r3/t2/t2/s0/out_reg_n_18 ,\r3/t2/t2/s0/out_reg_n_19 ,\r3/t2/t2/s0/out_reg_n_20 ,\r3/t2/t2/s0/out_reg_n_21 ,\r3/t2/t2/s0/out_reg_n_22 ,\r3/t2/t2/s0/out_reg_n_23 ,\r3/t2/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r3/t2/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[47:40],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[39:32],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r3/t2/t2/s4/out_reg_n_0 ,\r3/t2/t2/s4/out_reg_n_1 ,\r3/t2/t2/s4/out_reg_n_2 ,\r3/t2/t2/s4/out_reg_n_3 ,\r3/t2/t2/s4/out_reg_n_4 ,\r3/t2/t2/s4/out_reg_n_5 ,\r3/t2/t2/s4/out_reg_n_6 ,\r3/t2/t2/s4/out_reg_n_7 ,\r3/t2/t2/p_1_in }),
        .DOBDO({\r3/t2/t2/s4/out_reg_n_16 ,\r3/t2/t2/s4/out_reg_n_17 ,\r3/t2/t2/s4/out_reg_n_18 ,\r3/t2/t2/s4/out_reg_n_19 ,\r3/t2/t2/s4/out_reg_n_20 ,\r3/t2/t2/s4/out_reg_n_21 ,\r3/t2/t2/s4/out_reg_n_22 ,\r3/t2/t2/s4/out_reg_n_23 ,\r3/t2/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r3/t3/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r3/t3/t0/s0/out_reg_n_0 ,\r3/t3/t0/s0/out_reg_n_1 ,\r3/t3/t0/s0/out_reg_n_2 ,\r3/t3/t0/s0/out_reg_n_3 ,\r3/t3/t0/s0/out_reg_n_4 ,\r3/t3/t0/s0/out_reg_n_5 ,\r3/t3/t0/s0/out_reg_n_6 ,\r3/t3/t0/s0/out_reg_n_7 ,\r3/t3/t0/p_0_in }),
        .DOBDO({\r3/t3/t0/s0/out_reg_n_16 ,\r3/t3/t0/s0/out_reg_n_17 ,\r3/t3/t0/s0/out_reg_n_18 ,\r3/t3/t0/s0/out_reg_n_19 ,\r3/t3/t0/s0/out_reg_n_20 ,\r3/t3/t0/s0/out_reg_n_21 ,\r3/t3/t0/s0/out_reg_n_22 ,\r3/t3/t0/s0/out_reg_n_23 ,\r3/t3/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r3/t3/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r3/t3/t0/s4/out_reg_n_0 ,\r3/t3/t0/s4/out_reg_n_1 ,\r3/t3/t0/s4/out_reg_n_2 ,\r3/t3/t0/s4/out_reg_n_3 ,\r3/t3/t0/s4/out_reg_n_4 ,\r3/t3/t0/s4/out_reg_n_5 ,\r3/t3/t0/s4/out_reg_n_6 ,\r3/t3/t0/s4/out_reg_n_7 ,\r3/t3/t0/p_1_in }),
        .DOBDO({\r3/t3/t0/s4/out_reg_n_16 ,\r3/t3/t0/s4/out_reg_n_17 ,\r3/t3/t0/s4/out_reg_n_18 ,\r3/t3/t0/s4/out_reg_n_19 ,\r3/t3/t0/s4/out_reg_n_20 ,\r3/t3/t0/s4/out_reg_n_21 ,\r3/t3/t0/s4/out_reg_n_22 ,\r3/t3/t0/s4/out_reg_n_23 ,\r3/t3/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r3/t3/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r3/t3/t2/s0/out_reg_n_0 ,\r3/t3/t2/s0/out_reg_n_1 ,\r3/t3/t2/s0/out_reg_n_2 ,\r3/t3/t2/s0/out_reg_n_3 ,\r3/t3/t2/s0/out_reg_n_4 ,\r3/t3/t2/s0/out_reg_n_5 ,\r3/t3/t2/s0/out_reg_n_6 ,\r3/t3/t2/s0/out_reg_n_7 ,\r3/t3/t2/p_0_in }),
        .DOBDO({\r3/t3/t2/s0/out_reg_n_16 ,\r3/t3/t2/s0/out_reg_n_17 ,\r3/t3/t2/s0/out_reg_n_18 ,\r3/t3/t2/s0/out_reg_n_19 ,\r3/t3/t2/s0/out_reg_n_20 ,\r3/t3/t2/s0/out_reg_n_21 ,\r3/t3/t2/s0/out_reg_n_22 ,\r3/t3/t2/s0/out_reg_n_23 ,\r3/t3/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r3/t3/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s2[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r3/t3/t2/s4/out_reg_n_0 ,\r3/t3/t2/s4/out_reg_n_1 ,\r3/t3/t2/s4/out_reg_n_2 ,\r3/t3/t2/s4/out_reg_n_3 ,\r3/t3/t2/s4/out_reg_n_4 ,\r3/t3/t2/s4/out_reg_n_5 ,\r3/t3/t2/s4/out_reg_n_6 ,\r3/t3/t2/s4/out_reg_n_7 ,\r3/t3/t2/p_1_in }),
        .DOBDO({\r3/t3/t2/s4/out_reg_n_16 ,\r3/t3/t2/s4/out_reg_n_17 ,\r3/t3/t2/s4/out_reg_n_18 ,\r3/t3/t2/s4/out_reg_n_19 ,\r3/t3/t2/s4/out_reg_n_20 ,\r3/t3/t2/s4/out_reg_n_21 ,\r3/t3/t2/s4/out_reg_n_22 ,\r3/t3/t2/s4/out_reg_n_23 ,\r3/t3/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [0]),
        .Q(s4[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[100] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [100]),
        .Q(s4[100]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[101] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [101]),
        .Q(s4[101]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[102] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [102]),
        .Q(s4[102]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[103] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [103]),
        .Q(s4[103]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[104] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [104]),
        .Q(s4[104]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[105] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [105]),
        .Q(s4[105]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[106] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [106]),
        .Q(s4[106]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[107] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [107]),
        .Q(s4[107]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[108] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [108]),
        .Q(s4[108]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[109] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [109]),
        .Q(s4[109]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [10]),
        .Q(s4[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[110] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [110]),
        .Q(s4[110]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[111] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [111]),
        .Q(s4[111]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[112] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [112]),
        .Q(s4[112]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[113] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [113]),
        .Q(s4[113]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[114] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [114]),
        .Q(s4[114]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[115] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [115]),
        .Q(s4[115]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[116] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [116]),
        .Q(s4[116]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[117] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [117]),
        .Q(s4[117]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[118] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [118]),
        .Q(s4[118]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[119] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [119]),
        .Q(s4[119]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [11]),
        .Q(s4[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[120] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [120]),
        .Q(s4[120]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[121] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [121]),
        .Q(s4[121]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[122] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [122]),
        .Q(s4[122]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[123] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [123]),
        .Q(s4[123]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[124] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [124]),
        .Q(s4[124]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[125] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [125]),
        .Q(s4[125]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[126] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [126]),
        .Q(s4[126]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[127] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [127]),
        .Q(s4[127]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [12]),
        .Q(s4[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [13]),
        .Q(s4[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [14]),
        .Q(s4[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [15]),
        .Q(s4[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [16]),
        .Q(s4[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [17]),
        .Q(s4[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [18]),
        .Q(s4[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [19]),
        .Q(s4[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [1]),
        .Q(s4[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [20]),
        .Q(s4[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [21]),
        .Q(s4[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [22]),
        .Q(s4[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [23]),
        .Q(s4[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [24]),
        .Q(s4[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [25]),
        .Q(s4[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [26]),
        .Q(s4[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [27]),
        .Q(s4[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [28]),
        .Q(s4[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [29]),
        .Q(s4[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [2]),
        .Q(s4[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [30]),
        .Q(s4[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [31]),
        .Q(s4[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [32]),
        .Q(s4[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [33]),
        .Q(s4[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [34]),
        .Q(s4[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [35]),
        .Q(s4[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [36]),
        .Q(s4[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [37]),
        .Q(s4[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [38]),
        .Q(s4[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [39]),
        .Q(s4[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [3]),
        .Q(s4[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [40]),
        .Q(s4[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [41]),
        .Q(s4[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [42]),
        .Q(s4[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [43]),
        .Q(s4[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [44]),
        .Q(s4[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [45]),
        .Q(s4[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [46]),
        .Q(s4[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [47]),
        .Q(s4[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [48]),
        .Q(s4[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [49]),
        .Q(s4[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [4]),
        .Q(s4[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [50]),
        .Q(s4[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [51]),
        .Q(s4[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [52]),
        .Q(s4[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [53]),
        .Q(s4[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [54]),
        .Q(s4[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [55]),
        .Q(s4[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [56]),
        .Q(s4[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [57]),
        .Q(s4[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [58]),
        .Q(s4[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [59]),
        .Q(s4[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [5]),
        .Q(s4[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [60]),
        .Q(s4[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [61]),
        .Q(s4[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [62]),
        .Q(s4[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [63]),
        .Q(s4[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[64] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [64]),
        .Q(s4[64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[65] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [65]),
        .Q(s4[65]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[66] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [66]),
        .Q(s4[66]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[67] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [67]),
        .Q(s4[67]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[68] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [68]),
        .Q(s4[68]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[69] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [69]),
        .Q(s4[69]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [6]),
        .Q(s4[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[70] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [70]),
        .Q(s4[70]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[71] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [71]),
        .Q(s4[71]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[72] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [72]),
        .Q(s4[72]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[73] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [73]),
        .Q(s4[73]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[74] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [74]),
        .Q(s4[74]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[75] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [75]),
        .Q(s4[75]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[76] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [76]),
        .Q(s4[76]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[77] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [77]),
        .Q(s4[77]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[78] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [78]),
        .Q(s4[78]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[79] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [79]),
        .Q(s4[79]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [7]),
        .Q(s4[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[80] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [80]),
        .Q(s4[80]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[81] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [81]),
        .Q(s4[81]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[82] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [82]),
        .Q(s4[82]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[83] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [83]),
        .Q(s4[83]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[84] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [84]),
        .Q(s4[84]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[85] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [85]),
        .Q(s4[85]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[86] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [86]),
        .Q(s4[86]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[87] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [87]),
        .Q(s4[87]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[88] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [88]),
        .Q(s4[88]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[89] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [89]),
        .Q(s4[89]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [8]),
        .Q(s4[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[90] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [90]),
        .Q(s4[90]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[91] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [91]),
        .Q(s4[91]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[92] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [92]),
        .Q(s4[92]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[93] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [93]),
        .Q(s4[93]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[94] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [94]),
        .Q(s4[94]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[95] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [95]),
        .Q(s4[95]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[96] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [96]),
        .Q(s4[96]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[97] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [97]),
        .Q(s4[97]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[98] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [98]),
        .Q(s4[98]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[99] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [99]),
        .Q(s4[99]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r4/state_out_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r4/p_0_out [9]),
        .Q(s4[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r4/t0/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[127:120],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[119:112],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r4/t0/t0/s0/out_reg_n_0 ,\r4/t0/t0/s0/out_reg_n_1 ,\r4/t0/t0/s0/out_reg_n_2 ,\r4/t0/t0/s0/out_reg_n_3 ,\r4/t0/t0/s0/out_reg_n_4 ,\r4/t0/t0/s0/out_reg_n_5 ,\r4/t0/t0/s0/out_reg_n_6 ,\r4/t0/t0/s0/out_reg_n_7 ,\r4/t0/t0/p_0_in }),
        .DOBDO({\r4/t0/t0/s0/out_reg_n_16 ,\r4/t0/t0/s0/out_reg_n_17 ,\r4/t0/t0/s0/out_reg_n_18 ,\r4/t0/t0/s0/out_reg_n_19 ,\r4/t0/t0/s0/out_reg_n_20 ,\r4/t0/t0/s0/out_reg_n_21 ,\r4/t0/t0/s0/out_reg_n_22 ,\r4/t0/t0/s0/out_reg_n_23 ,\r4/t0/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r4/t0/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[127:120],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[119:112],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r4/t0/t0/s4/out_reg_n_0 ,\r4/t0/t0/s4/out_reg_n_1 ,\r4/t0/t0/s4/out_reg_n_2 ,\r4/t0/t0/s4/out_reg_n_3 ,\r4/t0/t0/s4/out_reg_n_4 ,\r4/t0/t0/s4/out_reg_n_5 ,\r4/t0/t0/s4/out_reg_n_6 ,\r4/t0/t0/s4/out_reg_n_7 ,\r4/t0/t0/p_1_in }),
        .DOBDO({\r4/t0/t0/s4/out_reg_n_16 ,\r4/t0/t0/s4/out_reg_n_17 ,\r4/t0/t0/s4/out_reg_n_18 ,\r4/t0/t0/s4/out_reg_n_19 ,\r4/t0/t0/s4/out_reg_n_20 ,\r4/t0/t0/s4/out_reg_n_21 ,\r4/t0/t0/s4/out_reg_n_22 ,\r4/t0/t0/s4/out_reg_n_23 ,\r4/t0/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r4/t0/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[111:104],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[103:96],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r4/t0/t2/s0/out_reg_n_0 ,\r4/t0/t2/s0/out_reg_n_1 ,\r4/t0/t2/s0/out_reg_n_2 ,\r4/t0/t2/s0/out_reg_n_3 ,\r4/t0/t2/s0/out_reg_n_4 ,\r4/t0/t2/s0/out_reg_n_5 ,\r4/t0/t2/s0/out_reg_n_6 ,\r4/t0/t2/s0/out_reg_n_7 ,\r4/t0/t2/p_0_in }),
        .DOBDO({\r4/t0/t2/s0/out_reg_n_16 ,\r4/t0/t2/s0/out_reg_n_17 ,\r4/t0/t2/s0/out_reg_n_18 ,\r4/t0/t2/s0/out_reg_n_19 ,\r4/t0/t2/s0/out_reg_n_20 ,\r4/t0/t2/s0/out_reg_n_21 ,\r4/t0/t2/s0/out_reg_n_22 ,\r4/t0/t2/s0/out_reg_n_23 ,\r4/t0/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r4/t0/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[111:104],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[103:96],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r4/t0/t2/s4/out_reg_n_0 ,\r4/t0/t2/s4/out_reg_n_1 ,\r4/t0/t2/s4/out_reg_n_2 ,\r4/t0/t2/s4/out_reg_n_3 ,\r4/t0/t2/s4/out_reg_n_4 ,\r4/t0/t2/s4/out_reg_n_5 ,\r4/t0/t2/s4/out_reg_n_6 ,\r4/t0/t2/s4/out_reg_n_7 ,\r4/t0/t2/p_1_in }),
        .DOBDO({\r4/t0/t2/s4/out_reg_n_16 ,\r4/t0/t2/s4/out_reg_n_17 ,\r4/t0/t2/s4/out_reg_n_18 ,\r4/t0/t2/s4/out_reg_n_19 ,\r4/t0/t2/s4/out_reg_n_20 ,\r4/t0/t2/s4/out_reg_n_21 ,\r4/t0/t2/s4/out_reg_n_22 ,\r4/t0/t2/s4/out_reg_n_23 ,\r4/t0/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r4/t1/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[95:88],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[87:80],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r4/t1/t0/s0/out_reg_n_0 ,\r4/t1/t0/s0/out_reg_n_1 ,\r4/t1/t0/s0/out_reg_n_2 ,\r4/t1/t0/s0/out_reg_n_3 ,\r4/t1/t0/s0/out_reg_n_4 ,\r4/t1/t0/s0/out_reg_n_5 ,\r4/t1/t0/s0/out_reg_n_6 ,\r4/t1/t0/s0/out_reg_n_7 ,\r4/t1/t0/p_0_in }),
        .DOBDO({\r4/t1/t0/s0/out_reg_n_16 ,\r4/t1/t0/s0/out_reg_n_17 ,\r4/t1/t0/s0/out_reg_n_18 ,\r4/t1/t0/s0/out_reg_n_19 ,\r4/t1/t0/s0/out_reg_n_20 ,\r4/t1/t0/s0/out_reg_n_21 ,\r4/t1/t0/s0/out_reg_n_22 ,\r4/t1/t0/s0/out_reg_n_23 ,\r4/t1/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r4/t1/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[95:88],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[87:80],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r4/t1/t0/s4/out_reg_n_0 ,\r4/t1/t0/s4/out_reg_n_1 ,\r4/t1/t0/s4/out_reg_n_2 ,\r4/t1/t0/s4/out_reg_n_3 ,\r4/t1/t0/s4/out_reg_n_4 ,\r4/t1/t0/s4/out_reg_n_5 ,\r4/t1/t0/s4/out_reg_n_6 ,\r4/t1/t0/s4/out_reg_n_7 ,\r4/t1/t0/p_1_in }),
        .DOBDO({\r4/t1/t0/s4/out_reg_n_16 ,\r4/t1/t0/s4/out_reg_n_17 ,\r4/t1/t0/s4/out_reg_n_18 ,\r4/t1/t0/s4/out_reg_n_19 ,\r4/t1/t0/s4/out_reg_n_20 ,\r4/t1/t0/s4/out_reg_n_21 ,\r4/t1/t0/s4/out_reg_n_22 ,\r4/t1/t0/s4/out_reg_n_23 ,\r4/t1/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r4/t1/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[79:72],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[71:64],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r4/t1/t2/s0/out_reg_n_0 ,\r4/t1/t2/s0/out_reg_n_1 ,\r4/t1/t2/s0/out_reg_n_2 ,\r4/t1/t2/s0/out_reg_n_3 ,\r4/t1/t2/s0/out_reg_n_4 ,\r4/t1/t2/s0/out_reg_n_5 ,\r4/t1/t2/s0/out_reg_n_6 ,\r4/t1/t2/s0/out_reg_n_7 ,\r4/t1/t2/p_0_in }),
        .DOBDO({\r4/t1/t2/s0/out_reg_n_16 ,\r4/t1/t2/s0/out_reg_n_17 ,\r4/t1/t2/s0/out_reg_n_18 ,\r4/t1/t2/s0/out_reg_n_19 ,\r4/t1/t2/s0/out_reg_n_20 ,\r4/t1/t2/s0/out_reg_n_21 ,\r4/t1/t2/s0/out_reg_n_22 ,\r4/t1/t2/s0/out_reg_n_23 ,\r4/t1/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r4/t1/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[79:72],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[71:64],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r4/t1/t2/s4/out_reg_n_0 ,\r4/t1/t2/s4/out_reg_n_1 ,\r4/t1/t2/s4/out_reg_n_2 ,\r4/t1/t2/s4/out_reg_n_3 ,\r4/t1/t2/s4/out_reg_n_4 ,\r4/t1/t2/s4/out_reg_n_5 ,\r4/t1/t2/s4/out_reg_n_6 ,\r4/t1/t2/s4/out_reg_n_7 ,\r4/t1/t2/p_1_in }),
        .DOBDO({\r4/t1/t2/s4/out_reg_n_16 ,\r4/t1/t2/s4/out_reg_n_17 ,\r4/t1/t2/s4/out_reg_n_18 ,\r4/t1/t2/s4/out_reg_n_19 ,\r4/t1/t2/s4/out_reg_n_20 ,\r4/t1/t2/s4/out_reg_n_21 ,\r4/t1/t2/s4/out_reg_n_22 ,\r4/t1/t2/s4/out_reg_n_23 ,\r4/t1/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r4/t2/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[63:56],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[55:48],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r4/t2/t0/s0/out_reg_n_0 ,\r4/t2/t0/s0/out_reg_n_1 ,\r4/t2/t0/s0/out_reg_n_2 ,\r4/t2/t0/s0/out_reg_n_3 ,\r4/t2/t0/s0/out_reg_n_4 ,\r4/t2/t0/s0/out_reg_n_5 ,\r4/t2/t0/s0/out_reg_n_6 ,\r4/t2/t0/s0/out_reg_n_7 ,\r4/t2/t0/p_0_in }),
        .DOBDO({\r4/t2/t0/s0/out_reg_n_16 ,\r4/t2/t0/s0/out_reg_n_17 ,\r4/t2/t0/s0/out_reg_n_18 ,\r4/t2/t0/s0/out_reg_n_19 ,\r4/t2/t0/s0/out_reg_n_20 ,\r4/t2/t0/s0/out_reg_n_21 ,\r4/t2/t0/s0/out_reg_n_22 ,\r4/t2/t0/s0/out_reg_n_23 ,\r4/t2/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r4/t2/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[63:56],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[55:48],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r4/t2/t0/s4/out_reg_n_0 ,\r4/t2/t0/s4/out_reg_n_1 ,\r4/t2/t0/s4/out_reg_n_2 ,\r4/t2/t0/s4/out_reg_n_3 ,\r4/t2/t0/s4/out_reg_n_4 ,\r4/t2/t0/s4/out_reg_n_5 ,\r4/t2/t0/s4/out_reg_n_6 ,\r4/t2/t0/s4/out_reg_n_7 ,\r4/t2/t0/p_1_in }),
        .DOBDO({\r4/t2/t0/s4/out_reg_n_16 ,\r4/t2/t0/s4/out_reg_n_17 ,\r4/t2/t0/s4/out_reg_n_18 ,\r4/t2/t0/s4/out_reg_n_19 ,\r4/t2/t0/s4/out_reg_n_20 ,\r4/t2/t0/s4/out_reg_n_21 ,\r4/t2/t0/s4/out_reg_n_22 ,\r4/t2/t0/s4/out_reg_n_23 ,\r4/t2/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r4/t2/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[47:40],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[39:32],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r4/t2/t2/s0/out_reg_n_0 ,\r4/t2/t2/s0/out_reg_n_1 ,\r4/t2/t2/s0/out_reg_n_2 ,\r4/t2/t2/s0/out_reg_n_3 ,\r4/t2/t2/s0/out_reg_n_4 ,\r4/t2/t2/s0/out_reg_n_5 ,\r4/t2/t2/s0/out_reg_n_6 ,\r4/t2/t2/s0/out_reg_n_7 ,\r4/t2/t2/p_0_in }),
        .DOBDO({\r4/t2/t2/s0/out_reg_n_16 ,\r4/t2/t2/s0/out_reg_n_17 ,\r4/t2/t2/s0/out_reg_n_18 ,\r4/t2/t2/s0/out_reg_n_19 ,\r4/t2/t2/s0/out_reg_n_20 ,\r4/t2/t2/s0/out_reg_n_21 ,\r4/t2/t2/s0/out_reg_n_22 ,\r4/t2/t2/s0/out_reg_n_23 ,\r4/t2/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r4/t2/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[47:40],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[39:32],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r4/t2/t2/s4/out_reg_n_0 ,\r4/t2/t2/s4/out_reg_n_1 ,\r4/t2/t2/s4/out_reg_n_2 ,\r4/t2/t2/s4/out_reg_n_3 ,\r4/t2/t2/s4/out_reg_n_4 ,\r4/t2/t2/s4/out_reg_n_5 ,\r4/t2/t2/s4/out_reg_n_6 ,\r4/t2/t2/s4/out_reg_n_7 ,\r4/t2/t2/p_1_in }),
        .DOBDO({\r4/t2/t2/s4/out_reg_n_16 ,\r4/t2/t2/s4/out_reg_n_17 ,\r4/t2/t2/s4/out_reg_n_18 ,\r4/t2/t2/s4/out_reg_n_19 ,\r4/t2/t2/s4/out_reg_n_20 ,\r4/t2/t2/s4/out_reg_n_21 ,\r4/t2/t2/s4/out_reg_n_22 ,\r4/t2/t2/s4/out_reg_n_23 ,\r4/t2/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r4/t3/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r4/t3/t0/s0/out_reg_n_0 ,\r4/t3/t0/s0/out_reg_n_1 ,\r4/t3/t0/s0/out_reg_n_2 ,\r4/t3/t0/s0/out_reg_n_3 ,\r4/t3/t0/s0/out_reg_n_4 ,\r4/t3/t0/s0/out_reg_n_5 ,\r4/t3/t0/s0/out_reg_n_6 ,\r4/t3/t0/s0/out_reg_n_7 ,\r4/t3/t0/p_0_in }),
        .DOBDO({\r4/t3/t0/s0/out_reg_n_16 ,\r4/t3/t0/s0/out_reg_n_17 ,\r4/t3/t0/s0/out_reg_n_18 ,\r4/t3/t0/s0/out_reg_n_19 ,\r4/t3/t0/s0/out_reg_n_20 ,\r4/t3/t0/s0/out_reg_n_21 ,\r4/t3/t0/s0/out_reg_n_22 ,\r4/t3/t0/s0/out_reg_n_23 ,\r4/t3/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r4/t3/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r4/t3/t0/s4/out_reg_n_0 ,\r4/t3/t0/s4/out_reg_n_1 ,\r4/t3/t0/s4/out_reg_n_2 ,\r4/t3/t0/s4/out_reg_n_3 ,\r4/t3/t0/s4/out_reg_n_4 ,\r4/t3/t0/s4/out_reg_n_5 ,\r4/t3/t0/s4/out_reg_n_6 ,\r4/t3/t0/s4/out_reg_n_7 ,\r4/t3/t0/p_1_in }),
        .DOBDO({\r4/t3/t0/s4/out_reg_n_16 ,\r4/t3/t0/s4/out_reg_n_17 ,\r4/t3/t0/s4/out_reg_n_18 ,\r4/t3/t0/s4/out_reg_n_19 ,\r4/t3/t0/s4/out_reg_n_20 ,\r4/t3/t0/s4/out_reg_n_21 ,\r4/t3/t0/s4/out_reg_n_22 ,\r4/t3/t0/s4/out_reg_n_23 ,\r4/t3/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r4/t3/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r4/t3/t2/s0/out_reg_n_0 ,\r4/t3/t2/s0/out_reg_n_1 ,\r4/t3/t2/s0/out_reg_n_2 ,\r4/t3/t2/s0/out_reg_n_3 ,\r4/t3/t2/s0/out_reg_n_4 ,\r4/t3/t2/s0/out_reg_n_5 ,\r4/t3/t2/s0/out_reg_n_6 ,\r4/t3/t2/s0/out_reg_n_7 ,\r4/t3/t2/p_0_in }),
        .DOBDO({\r4/t3/t2/s0/out_reg_n_16 ,\r4/t3/t2/s0/out_reg_n_17 ,\r4/t3/t2/s0/out_reg_n_18 ,\r4/t3/t2/s0/out_reg_n_19 ,\r4/t3/t2/s0/out_reg_n_20 ,\r4/t3/t2/s0/out_reg_n_21 ,\r4/t3/t2/s0/out_reg_n_22 ,\r4/t3/t2/s0/out_reg_n_23 ,\r4/t3/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r4/t3/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s3[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r4/t3/t2/s4/out_reg_n_0 ,\r4/t3/t2/s4/out_reg_n_1 ,\r4/t3/t2/s4/out_reg_n_2 ,\r4/t3/t2/s4/out_reg_n_3 ,\r4/t3/t2/s4/out_reg_n_4 ,\r4/t3/t2/s4/out_reg_n_5 ,\r4/t3/t2/s4/out_reg_n_6 ,\r4/t3/t2/s4/out_reg_n_7 ,\r4/t3/t2/p_1_in }),
        .DOBDO({\r4/t3/t2/s4/out_reg_n_16 ,\r4/t3/t2/s4/out_reg_n_17 ,\r4/t3/t2/s4/out_reg_n_18 ,\r4/t3/t2/s4/out_reg_n_19 ,\r4/t3/t2/s4/out_reg_n_20 ,\r4/t3/t2/s4/out_reg_n_21 ,\r4/t3/t2/s4/out_reg_n_22 ,\r4/t3/t2/s4/out_reg_n_23 ,\r4/t3/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [0]),
        .Q(s5[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[100] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [100]),
        .Q(s5[100]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[101] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [101]),
        .Q(s5[101]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[102] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [102]),
        .Q(s5[102]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[103] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [103]),
        .Q(s5[103]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[104] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [104]),
        .Q(s5[104]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[105] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [105]),
        .Q(s5[105]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[106] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [106]),
        .Q(s5[106]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[107] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [107]),
        .Q(s5[107]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[108] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [108]),
        .Q(s5[108]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[109] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [109]),
        .Q(s5[109]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [10]),
        .Q(s5[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[110] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [110]),
        .Q(s5[110]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[111] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [111]),
        .Q(s5[111]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[112] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [112]),
        .Q(s5[112]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[113] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [113]),
        .Q(s5[113]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[114] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [114]),
        .Q(s5[114]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[115] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [115]),
        .Q(s5[115]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[116] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [116]),
        .Q(s5[116]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[117] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [117]),
        .Q(s5[117]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[118] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [118]),
        .Q(s5[118]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[119] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [119]),
        .Q(s5[119]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [11]),
        .Q(s5[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[120] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [120]),
        .Q(s5[120]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[121] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [121]),
        .Q(s5[121]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[122] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [122]),
        .Q(s5[122]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[123] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [123]),
        .Q(s5[123]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[124] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [124]),
        .Q(s5[124]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[125] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [125]),
        .Q(s5[125]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[126] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [126]),
        .Q(s5[126]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[127] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [127]),
        .Q(s5[127]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [12]),
        .Q(s5[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [13]),
        .Q(s5[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [14]),
        .Q(s5[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [15]),
        .Q(s5[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [16]),
        .Q(s5[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [17]),
        .Q(s5[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [18]),
        .Q(s5[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [19]),
        .Q(s5[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [1]),
        .Q(s5[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [20]),
        .Q(s5[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [21]),
        .Q(s5[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [22]),
        .Q(s5[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [23]),
        .Q(s5[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [24]),
        .Q(s5[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [25]),
        .Q(s5[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [26]),
        .Q(s5[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [27]),
        .Q(s5[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [28]),
        .Q(s5[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [29]),
        .Q(s5[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [2]),
        .Q(s5[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [30]),
        .Q(s5[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [31]),
        .Q(s5[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [32]),
        .Q(s5[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [33]),
        .Q(s5[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [34]),
        .Q(s5[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [35]),
        .Q(s5[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [36]),
        .Q(s5[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [37]),
        .Q(s5[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [38]),
        .Q(s5[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [39]),
        .Q(s5[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [3]),
        .Q(s5[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [40]),
        .Q(s5[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [41]),
        .Q(s5[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [42]),
        .Q(s5[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [43]),
        .Q(s5[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [44]),
        .Q(s5[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [45]),
        .Q(s5[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [46]),
        .Q(s5[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [47]),
        .Q(s5[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [48]),
        .Q(s5[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [49]),
        .Q(s5[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [4]),
        .Q(s5[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [50]),
        .Q(s5[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [51]),
        .Q(s5[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [52]),
        .Q(s5[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [53]),
        .Q(s5[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [54]),
        .Q(s5[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [55]),
        .Q(s5[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [56]),
        .Q(s5[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [57]),
        .Q(s5[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [58]),
        .Q(s5[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [59]),
        .Q(s5[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [5]),
        .Q(s5[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [60]),
        .Q(s5[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [61]),
        .Q(s5[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [62]),
        .Q(s5[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [63]),
        .Q(s5[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[64] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [64]),
        .Q(s5[64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[65] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [65]),
        .Q(s5[65]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[66] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [66]),
        .Q(s5[66]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[67] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [67]),
        .Q(s5[67]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[68] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [68]),
        .Q(s5[68]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[69] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [69]),
        .Q(s5[69]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [6]),
        .Q(s5[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[70] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [70]),
        .Q(s5[70]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[71] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [71]),
        .Q(s5[71]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[72] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [72]),
        .Q(s5[72]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[73] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [73]),
        .Q(s5[73]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[74] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [74]),
        .Q(s5[74]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[75] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [75]),
        .Q(s5[75]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[76] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [76]),
        .Q(s5[76]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[77] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [77]),
        .Q(s5[77]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[78] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [78]),
        .Q(s5[78]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[79] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [79]),
        .Q(s5[79]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [7]),
        .Q(s5[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[80] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [80]),
        .Q(s5[80]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[81] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [81]),
        .Q(s5[81]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[82] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [82]),
        .Q(s5[82]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[83] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [83]),
        .Q(s5[83]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[84] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [84]),
        .Q(s5[84]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[85] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [85]),
        .Q(s5[85]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[86] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [86]),
        .Q(s5[86]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[87] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [87]),
        .Q(s5[87]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[88] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [88]),
        .Q(s5[88]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[89] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [89]),
        .Q(s5[89]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [8]),
        .Q(s5[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[90] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [90]),
        .Q(s5[90]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[91] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [91]),
        .Q(s5[91]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[92] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [92]),
        .Q(s5[92]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[93] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [93]),
        .Q(s5[93]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[94] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [94]),
        .Q(s5[94]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[95] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [95]),
        .Q(s5[95]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[96] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [96]),
        .Q(s5[96]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[97] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [97]),
        .Q(s5[97]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[98] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [98]),
        .Q(s5[98]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[99] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [99]),
        .Q(s5[99]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r5/state_out_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r5/p_0_out [9]),
        .Q(s5[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r5/t0/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[127:120],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[119:112],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r5/t0/t0/s0/out_reg_n_0 ,\r5/t0/t0/s0/out_reg_n_1 ,\r5/t0/t0/s0/out_reg_n_2 ,\r5/t0/t0/s0/out_reg_n_3 ,\r5/t0/t0/s0/out_reg_n_4 ,\r5/t0/t0/s0/out_reg_n_5 ,\r5/t0/t0/s0/out_reg_n_6 ,\r5/t0/t0/s0/out_reg_n_7 ,\r5/t0/t0/p_0_in }),
        .DOBDO({\r5/t0/t0/s0/out_reg_n_16 ,\r5/t0/t0/s0/out_reg_n_17 ,\r5/t0/t0/s0/out_reg_n_18 ,\r5/t0/t0/s0/out_reg_n_19 ,\r5/t0/t0/s0/out_reg_n_20 ,\r5/t0/t0/s0/out_reg_n_21 ,\r5/t0/t0/s0/out_reg_n_22 ,\r5/t0/t0/s0/out_reg_n_23 ,\r5/t0/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r5/t0/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[127:120],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[119:112],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r5/t0/t0/s4/out_reg_n_0 ,\r5/t0/t0/s4/out_reg_n_1 ,\r5/t0/t0/s4/out_reg_n_2 ,\r5/t0/t0/s4/out_reg_n_3 ,\r5/t0/t0/s4/out_reg_n_4 ,\r5/t0/t0/s4/out_reg_n_5 ,\r5/t0/t0/s4/out_reg_n_6 ,\r5/t0/t0/s4/out_reg_n_7 ,\r5/t0/t0/p_1_in }),
        .DOBDO({\r5/t0/t0/s4/out_reg_n_16 ,\r5/t0/t0/s4/out_reg_n_17 ,\r5/t0/t0/s4/out_reg_n_18 ,\r5/t0/t0/s4/out_reg_n_19 ,\r5/t0/t0/s4/out_reg_n_20 ,\r5/t0/t0/s4/out_reg_n_21 ,\r5/t0/t0/s4/out_reg_n_22 ,\r5/t0/t0/s4/out_reg_n_23 ,\r5/t0/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r5/t0/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[111:104],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[103:96],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r5/t0/t2/s0/out_reg_n_0 ,\r5/t0/t2/s0/out_reg_n_1 ,\r5/t0/t2/s0/out_reg_n_2 ,\r5/t0/t2/s0/out_reg_n_3 ,\r5/t0/t2/s0/out_reg_n_4 ,\r5/t0/t2/s0/out_reg_n_5 ,\r5/t0/t2/s0/out_reg_n_6 ,\r5/t0/t2/s0/out_reg_n_7 ,\r5/t0/t2/p_0_in }),
        .DOBDO({\r5/t0/t2/s0/out_reg_n_16 ,\r5/t0/t2/s0/out_reg_n_17 ,\r5/t0/t2/s0/out_reg_n_18 ,\r5/t0/t2/s0/out_reg_n_19 ,\r5/t0/t2/s0/out_reg_n_20 ,\r5/t0/t2/s0/out_reg_n_21 ,\r5/t0/t2/s0/out_reg_n_22 ,\r5/t0/t2/s0/out_reg_n_23 ,\r5/t0/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r5/t0/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[111:104],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[103:96],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r5/t0/t2/s4/out_reg_n_0 ,\r5/t0/t2/s4/out_reg_n_1 ,\r5/t0/t2/s4/out_reg_n_2 ,\r5/t0/t2/s4/out_reg_n_3 ,\r5/t0/t2/s4/out_reg_n_4 ,\r5/t0/t2/s4/out_reg_n_5 ,\r5/t0/t2/s4/out_reg_n_6 ,\r5/t0/t2/s4/out_reg_n_7 ,\r5/t0/t2/p_1_in }),
        .DOBDO({\r5/t0/t2/s4/out_reg_n_16 ,\r5/t0/t2/s4/out_reg_n_17 ,\r5/t0/t2/s4/out_reg_n_18 ,\r5/t0/t2/s4/out_reg_n_19 ,\r5/t0/t2/s4/out_reg_n_20 ,\r5/t0/t2/s4/out_reg_n_21 ,\r5/t0/t2/s4/out_reg_n_22 ,\r5/t0/t2/s4/out_reg_n_23 ,\r5/t0/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r5/t1/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[95:88],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[87:80],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r5/t1/t0/s0/out_reg_n_0 ,\r5/t1/t0/s0/out_reg_n_1 ,\r5/t1/t0/s0/out_reg_n_2 ,\r5/t1/t0/s0/out_reg_n_3 ,\r5/t1/t0/s0/out_reg_n_4 ,\r5/t1/t0/s0/out_reg_n_5 ,\r5/t1/t0/s0/out_reg_n_6 ,\r5/t1/t0/s0/out_reg_n_7 ,\r5/t1/t0/p_0_in }),
        .DOBDO({\r5/t1/t0/s0/out_reg_n_16 ,\r5/t1/t0/s0/out_reg_n_17 ,\r5/t1/t0/s0/out_reg_n_18 ,\r5/t1/t0/s0/out_reg_n_19 ,\r5/t1/t0/s0/out_reg_n_20 ,\r5/t1/t0/s0/out_reg_n_21 ,\r5/t1/t0/s0/out_reg_n_22 ,\r5/t1/t0/s0/out_reg_n_23 ,\r5/t1/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r5/t1/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[95:88],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[87:80],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r5/t1/t0/s4/out_reg_n_0 ,\r5/t1/t0/s4/out_reg_n_1 ,\r5/t1/t0/s4/out_reg_n_2 ,\r5/t1/t0/s4/out_reg_n_3 ,\r5/t1/t0/s4/out_reg_n_4 ,\r5/t1/t0/s4/out_reg_n_5 ,\r5/t1/t0/s4/out_reg_n_6 ,\r5/t1/t0/s4/out_reg_n_7 ,\r5/t1/t0/p_1_in }),
        .DOBDO({\r5/t1/t0/s4/out_reg_n_16 ,\r5/t1/t0/s4/out_reg_n_17 ,\r5/t1/t0/s4/out_reg_n_18 ,\r5/t1/t0/s4/out_reg_n_19 ,\r5/t1/t0/s4/out_reg_n_20 ,\r5/t1/t0/s4/out_reg_n_21 ,\r5/t1/t0/s4/out_reg_n_22 ,\r5/t1/t0/s4/out_reg_n_23 ,\r5/t1/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r5/t1/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[79:72],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[71:64],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r5/t1/t2/s0/out_reg_n_0 ,\r5/t1/t2/s0/out_reg_n_1 ,\r5/t1/t2/s0/out_reg_n_2 ,\r5/t1/t2/s0/out_reg_n_3 ,\r5/t1/t2/s0/out_reg_n_4 ,\r5/t1/t2/s0/out_reg_n_5 ,\r5/t1/t2/s0/out_reg_n_6 ,\r5/t1/t2/s0/out_reg_n_7 ,\r5/t1/t2/p_0_in }),
        .DOBDO({\r5/t1/t2/s0/out_reg_n_16 ,\r5/t1/t2/s0/out_reg_n_17 ,\r5/t1/t2/s0/out_reg_n_18 ,\r5/t1/t2/s0/out_reg_n_19 ,\r5/t1/t2/s0/out_reg_n_20 ,\r5/t1/t2/s0/out_reg_n_21 ,\r5/t1/t2/s0/out_reg_n_22 ,\r5/t1/t2/s0/out_reg_n_23 ,\r5/t1/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r5/t1/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[79:72],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[71:64],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r5/t1/t2/s4/out_reg_n_0 ,\r5/t1/t2/s4/out_reg_n_1 ,\r5/t1/t2/s4/out_reg_n_2 ,\r5/t1/t2/s4/out_reg_n_3 ,\r5/t1/t2/s4/out_reg_n_4 ,\r5/t1/t2/s4/out_reg_n_5 ,\r5/t1/t2/s4/out_reg_n_6 ,\r5/t1/t2/s4/out_reg_n_7 ,\r5/t1/t2/p_1_in }),
        .DOBDO({\r5/t1/t2/s4/out_reg_n_16 ,\r5/t1/t2/s4/out_reg_n_17 ,\r5/t1/t2/s4/out_reg_n_18 ,\r5/t1/t2/s4/out_reg_n_19 ,\r5/t1/t2/s4/out_reg_n_20 ,\r5/t1/t2/s4/out_reg_n_21 ,\r5/t1/t2/s4/out_reg_n_22 ,\r5/t1/t2/s4/out_reg_n_23 ,\r5/t1/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r5/t2/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[63:56],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[55:48],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r5/t2/t0/s0/out_reg_n_0 ,\r5/t2/t0/s0/out_reg_n_1 ,\r5/t2/t0/s0/out_reg_n_2 ,\r5/t2/t0/s0/out_reg_n_3 ,\r5/t2/t0/s0/out_reg_n_4 ,\r5/t2/t0/s0/out_reg_n_5 ,\r5/t2/t0/s0/out_reg_n_6 ,\r5/t2/t0/s0/out_reg_n_7 ,\r5/t2/t0/p_0_in }),
        .DOBDO({\r5/t2/t0/s0/out_reg_n_16 ,\r5/t2/t0/s0/out_reg_n_17 ,\r5/t2/t0/s0/out_reg_n_18 ,\r5/t2/t0/s0/out_reg_n_19 ,\r5/t2/t0/s0/out_reg_n_20 ,\r5/t2/t0/s0/out_reg_n_21 ,\r5/t2/t0/s0/out_reg_n_22 ,\r5/t2/t0/s0/out_reg_n_23 ,\r5/t2/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r5/t2/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[63:56],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[55:48],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r5/t2/t0/s4/out_reg_n_0 ,\r5/t2/t0/s4/out_reg_n_1 ,\r5/t2/t0/s4/out_reg_n_2 ,\r5/t2/t0/s4/out_reg_n_3 ,\r5/t2/t0/s4/out_reg_n_4 ,\r5/t2/t0/s4/out_reg_n_5 ,\r5/t2/t0/s4/out_reg_n_6 ,\r5/t2/t0/s4/out_reg_n_7 ,\r5/t2/t0/p_1_in }),
        .DOBDO({\r5/t2/t0/s4/out_reg_n_16 ,\r5/t2/t0/s4/out_reg_n_17 ,\r5/t2/t0/s4/out_reg_n_18 ,\r5/t2/t0/s4/out_reg_n_19 ,\r5/t2/t0/s4/out_reg_n_20 ,\r5/t2/t0/s4/out_reg_n_21 ,\r5/t2/t0/s4/out_reg_n_22 ,\r5/t2/t0/s4/out_reg_n_23 ,\r5/t2/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r5/t2/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[47:40],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[39:32],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r5/t2/t2/s0/out_reg_n_0 ,\r5/t2/t2/s0/out_reg_n_1 ,\r5/t2/t2/s0/out_reg_n_2 ,\r5/t2/t2/s0/out_reg_n_3 ,\r5/t2/t2/s0/out_reg_n_4 ,\r5/t2/t2/s0/out_reg_n_5 ,\r5/t2/t2/s0/out_reg_n_6 ,\r5/t2/t2/s0/out_reg_n_7 ,\r5/t2/t2/p_0_in }),
        .DOBDO({\r5/t2/t2/s0/out_reg_n_16 ,\r5/t2/t2/s0/out_reg_n_17 ,\r5/t2/t2/s0/out_reg_n_18 ,\r5/t2/t2/s0/out_reg_n_19 ,\r5/t2/t2/s0/out_reg_n_20 ,\r5/t2/t2/s0/out_reg_n_21 ,\r5/t2/t2/s0/out_reg_n_22 ,\r5/t2/t2/s0/out_reg_n_23 ,\r5/t2/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r5/t2/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[47:40],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[39:32],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r5/t2/t2/s4/out_reg_n_0 ,\r5/t2/t2/s4/out_reg_n_1 ,\r5/t2/t2/s4/out_reg_n_2 ,\r5/t2/t2/s4/out_reg_n_3 ,\r5/t2/t2/s4/out_reg_n_4 ,\r5/t2/t2/s4/out_reg_n_5 ,\r5/t2/t2/s4/out_reg_n_6 ,\r5/t2/t2/s4/out_reg_n_7 ,\r5/t2/t2/p_1_in }),
        .DOBDO({\r5/t2/t2/s4/out_reg_n_16 ,\r5/t2/t2/s4/out_reg_n_17 ,\r5/t2/t2/s4/out_reg_n_18 ,\r5/t2/t2/s4/out_reg_n_19 ,\r5/t2/t2/s4/out_reg_n_20 ,\r5/t2/t2/s4/out_reg_n_21 ,\r5/t2/t2/s4/out_reg_n_22 ,\r5/t2/t2/s4/out_reg_n_23 ,\r5/t2/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r5/t3/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r5/t3/t0/s0/out_reg_n_0 ,\r5/t3/t0/s0/out_reg_n_1 ,\r5/t3/t0/s0/out_reg_n_2 ,\r5/t3/t0/s0/out_reg_n_3 ,\r5/t3/t0/s0/out_reg_n_4 ,\r5/t3/t0/s0/out_reg_n_5 ,\r5/t3/t0/s0/out_reg_n_6 ,\r5/t3/t0/s0/out_reg_n_7 ,\r5/t3/t0/p_0_in }),
        .DOBDO({\r5/t3/t0/s0/out_reg_n_16 ,\r5/t3/t0/s0/out_reg_n_17 ,\r5/t3/t0/s0/out_reg_n_18 ,\r5/t3/t0/s0/out_reg_n_19 ,\r5/t3/t0/s0/out_reg_n_20 ,\r5/t3/t0/s0/out_reg_n_21 ,\r5/t3/t0/s0/out_reg_n_22 ,\r5/t3/t0/s0/out_reg_n_23 ,\r5/t3/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r5/t3/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r5/t3/t0/s4/out_reg_n_0 ,\r5/t3/t0/s4/out_reg_n_1 ,\r5/t3/t0/s4/out_reg_n_2 ,\r5/t3/t0/s4/out_reg_n_3 ,\r5/t3/t0/s4/out_reg_n_4 ,\r5/t3/t0/s4/out_reg_n_5 ,\r5/t3/t0/s4/out_reg_n_6 ,\r5/t3/t0/s4/out_reg_n_7 ,\r5/t3/t0/p_1_in }),
        .DOBDO({\r5/t3/t0/s4/out_reg_n_16 ,\r5/t3/t0/s4/out_reg_n_17 ,\r5/t3/t0/s4/out_reg_n_18 ,\r5/t3/t0/s4/out_reg_n_19 ,\r5/t3/t0/s4/out_reg_n_20 ,\r5/t3/t0/s4/out_reg_n_21 ,\r5/t3/t0/s4/out_reg_n_22 ,\r5/t3/t0/s4/out_reg_n_23 ,\r5/t3/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r5/t3/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r5/t3/t2/s0/out_reg_n_0 ,\r5/t3/t2/s0/out_reg_n_1 ,\r5/t3/t2/s0/out_reg_n_2 ,\r5/t3/t2/s0/out_reg_n_3 ,\r5/t3/t2/s0/out_reg_n_4 ,\r5/t3/t2/s0/out_reg_n_5 ,\r5/t3/t2/s0/out_reg_n_6 ,\r5/t3/t2/s0/out_reg_n_7 ,\r5/t3/t2/p_0_in }),
        .DOBDO({\r5/t3/t2/s0/out_reg_n_16 ,\r5/t3/t2/s0/out_reg_n_17 ,\r5/t3/t2/s0/out_reg_n_18 ,\r5/t3/t2/s0/out_reg_n_19 ,\r5/t3/t2/s0/out_reg_n_20 ,\r5/t3/t2/s0/out_reg_n_21 ,\r5/t3/t2/s0/out_reg_n_22 ,\r5/t3/t2/s0/out_reg_n_23 ,\r5/t3/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r5/t3/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s4[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r5/t3/t2/s4/out_reg_n_0 ,\r5/t3/t2/s4/out_reg_n_1 ,\r5/t3/t2/s4/out_reg_n_2 ,\r5/t3/t2/s4/out_reg_n_3 ,\r5/t3/t2/s4/out_reg_n_4 ,\r5/t3/t2/s4/out_reg_n_5 ,\r5/t3/t2/s4/out_reg_n_6 ,\r5/t3/t2/s4/out_reg_n_7 ,\r5/t3/t2/p_1_in }),
        .DOBDO({\r5/t3/t2/s4/out_reg_n_16 ,\r5/t3/t2/s4/out_reg_n_17 ,\r5/t3/t2/s4/out_reg_n_18 ,\r5/t3/t2/s4/out_reg_n_19 ,\r5/t3/t2/s4/out_reg_n_20 ,\r5/t3/t2/s4/out_reg_n_21 ,\r5/t3/t2/s4/out_reg_n_22 ,\r5/t3/t2/s4/out_reg_n_23 ,\r5/t3/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [0]),
        .Q(s6[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[100] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [100]),
        .Q(s6[100]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[101] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [101]),
        .Q(s6[101]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[102] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [102]),
        .Q(s6[102]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[103] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [103]),
        .Q(s6[103]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[104] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [104]),
        .Q(s6[104]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[105] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [105]),
        .Q(s6[105]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[106] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [106]),
        .Q(s6[106]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[107] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [107]),
        .Q(s6[107]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[108] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [108]),
        .Q(s6[108]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[109] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [109]),
        .Q(s6[109]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [10]),
        .Q(s6[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[110] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [110]),
        .Q(s6[110]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[111] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [111]),
        .Q(s6[111]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[112] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [112]),
        .Q(s6[112]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[113] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [113]),
        .Q(s6[113]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[114] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [114]),
        .Q(s6[114]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[115] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [115]),
        .Q(s6[115]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[116] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [116]),
        .Q(s6[116]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[117] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [117]),
        .Q(s6[117]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[118] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [118]),
        .Q(s6[118]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[119] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [119]),
        .Q(s6[119]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [11]),
        .Q(s6[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[120] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [120]),
        .Q(s6[120]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[121] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [121]),
        .Q(s6[121]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[122] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [122]),
        .Q(s6[122]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[123] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [123]),
        .Q(s6[123]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[124] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [124]),
        .Q(s6[124]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[125] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [125]),
        .Q(s6[125]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[126] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [126]),
        .Q(s6[126]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[127] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [127]),
        .Q(s6[127]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [12]),
        .Q(s6[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [13]),
        .Q(s6[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [14]),
        .Q(s6[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [15]),
        .Q(s6[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [16]),
        .Q(s6[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [17]),
        .Q(s6[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [18]),
        .Q(s6[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [19]),
        .Q(s6[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [1]),
        .Q(s6[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [20]),
        .Q(s6[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [21]),
        .Q(s6[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [22]),
        .Q(s6[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [23]),
        .Q(s6[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [24]),
        .Q(s6[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [25]),
        .Q(s6[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [26]),
        .Q(s6[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [27]),
        .Q(s6[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [28]),
        .Q(s6[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [29]),
        .Q(s6[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [2]),
        .Q(s6[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [30]),
        .Q(s6[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [31]),
        .Q(s6[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [32]),
        .Q(s6[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [33]),
        .Q(s6[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [34]),
        .Q(s6[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [35]),
        .Q(s6[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [36]),
        .Q(s6[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [37]),
        .Q(s6[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [38]),
        .Q(s6[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [39]),
        .Q(s6[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [3]),
        .Q(s6[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [40]),
        .Q(s6[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [41]),
        .Q(s6[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [42]),
        .Q(s6[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [43]),
        .Q(s6[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [44]),
        .Q(s6[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [45]),
        .Q(s6[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [46]),
        .Q(s6[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [47]),
        .Q(s6[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [48]),
        .Q(s6[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [49]),
        .Q(s6[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [4]),
        .Q(s6[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [50]),
        .Q(s6[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [51]),
        .Q(s6[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [52]),
        .Q(s6[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [53]),
        .Q(s6[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [54]),
        .Q(s6[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [55]),
        .Q(s6[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [56]),
        .Q(s6[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [57]),
        .Q(s6[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [58]),
        .Q(s6[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [59]),
        .Q(s6[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [5]),
        .Q(s6[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [60]),
        .Q(s6[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [61]),
        .Q(s6[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [62]),
        .Q(s6[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [63]),
        .Q(s6[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[64] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [64]),
        .Q(s6[64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[65] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [65]),
        .Q(s6[65]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[66] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [66]),
        .Q(s6[66]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[67] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [67]),
        .Q(s6[67]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[68] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [68]),
        .Q(s6[68]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[69] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [69]),
        .Q(s6[69]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [6]),
        .Q(s6[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[70] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [70]),
        .Q(s6[70]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[71] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [71]),
        .Q(s6[71]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[72] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [72]),
        .Q(s6[72]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[73] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [73]),
        .Q(s6[73]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[74] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [74]),
        .Q(s6[74]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[75] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [75]),
        .Q(s6[75]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[76] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [76]),
        .Q(s6[76]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[77] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [77]),
        .Q(s6[77]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[78] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [78]),
        .Q(s6[78]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[79] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [79]),
        .Q(s6[79]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [7]),
        .Q(s6[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[80] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [80]),
        .Q(s6[80]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[81] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [81]),
        .Q(s6[81]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[82] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [82]),
        .Q(s6[82]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[83] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [83]),
        .Q(s6[83]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[84] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [84]),
        .Q(s6[84]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[85] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [85]),
        .Q(s6[85]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[86] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [86]),
        .Q(s6[86]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[87] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [87]),
        .Q(s6[87]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[88] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [88]),
        .Q(s6[88]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[89] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [89]),
        .Q(s6[89]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [8]),
        .Q(s6[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[90] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [90]),
        .Q(s6[90]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[91] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [91]),
        .Q(s6[91]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[92] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [92]),
        .Q(s6[92]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[93] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [93]),
        .Q(s6[93]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[94] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [94]),
        .Q(s6[94]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[95] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [95]),
        .Q(s6[95]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[96] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [96]),
        .Q(s6[96]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[97] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [97]),
        .Q(s6[97]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[98] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [98]),
        .Q(s6[98]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[99] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [99]),
        .Q(s6[99]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r6/state_out_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r6/p_0_out [9]),
        .Q(s6[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r6/t0/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[127:120],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[119:112],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r6/t0/t0/s0/out_reg_n_0 ,\r6/t0/t0/s0/out_reg_n_1 ,\r6/t0/t0/s0/out_reg_n_2 ,\r6/t0/t0/s0/out_reg_n_3 ,\r6/t0/t0/s0/out_reg_n_4 ,\r6/t0/t0/s0/out_reg_n_5 ,\r6/t0/t0/s0/out_reg_n_6 ,\r6/t0/t0/s0/out_reg_n_7 ,\r6/t0/t0/p_0_in }),
        .DOBDO({\r6/t0/t0/s0/out_reg_n_16 ,\r6/t0/t0/s0/out_reg_n_17 ,\r6/t0/t0/s0/out_reg_n_18 ,\r6/t0/t0/s0/out_reg_n_19 ,\r6/t0/t0/s0/out_reg_n_20 ,\r6/t0/t0/s0/out_reg_n_21 ,\r6/t0/t0/s0/out_reg_n_22 ,\r6/t0/t0/s0/out_reg_n_23 ,\r6/t0/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r6/t0/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[127:120],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[119:112],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r6/t0/t0/s4/out_reg_n_0 ,\r6/t0/t0/s4/out_reg_n_1 ,\r6/t0/t0/s4/out_reg_n_2 ,\r6/t0/t0/s4/out_reg_n_3 ,\r6/t0/t0/s4/out_reg_n_4 ,\r6/t0/t0/s4/out_reg_n_5 ,\r6/t0/t0/s4/out_reg_n_6 ,\r6/t0/t0/s4/out_reg_n_7 ,\r6/t0/t0/p_1_in }),
        .DOBDO({\r6/t0/t0/s4/out_reg_n_16 ,\r6/t0/t0/s4/out_reg_n_17 ,\r6/t0/t0/s4/out_reg_n_18 ,\r6/t0/t0/s4/out_reg_n_19 ,\r6/t0/t0/s4/out_reg_n_20 ,\r6/t0/t0/s4/out_reg_n_21 ,\r6/t0/t0/s4/out_reg_n_22 ,\r6/t0/t0/s4/out_reg_n_23 ,\r6/t0/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r6/t0/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[111:104],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[103:96],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r6/t0/t2/s0/out_reg_n_0 ,\r6/t0/t2/s0/out_reg_n_1 ,\r6/t0/t2/s0/out_reg_n_2 ,\r6/t0/t2/s0/out_reg_n_3 ,\r6/t0/t2/s0/out_reg_n_4 ,\r6/t0/t2/s0/out_reg_n_5 ,\r6/t0/t2/s0/out_reg_n_6 ,\r6/t0/t2/s0/out_reg_n_7 ,\r6/t0/t2/p_0_in }),
        .DOBDO({\r6/t0/t2/s0/out_reg_n_16 ,\r6/t0/t2/s0/out_reg_n_17 ,\r6/t0/t2/s0/out_reg_n_18 ,\r6/t0/t2/s0/out_reg_n_19 ,\r6/t0/t2/s0/out_reg_n_20 ,\r6/t0/t2/s0/out_reg_n_21 ,\r6/t0/t2/s0/out_reg_n_22 ,\r6/t0/t2/s0/out_reg_n_23 ,\r6/t0/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r6/t0/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[111:104],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[103:96],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r6/t0/t2/s4/out_reg_n_0 ,\r6/t0/t2/s4/out_reg_n_1 ,\r6/t0/t2/s4/out_reg_n_2 ,\r6/t0/t2/s4/out_reg_n_3 ,\r6/t0/t2/s4/out_reg_n_4 ,\r6/t0/t2/s4/out_reg_n_5 ,\r6/t0/t2/s4/out_reg_n_6 ,\r6/t0/t2/s4/out_reg_n_7 ,\r6/t0/t2/p_1_in }),
        .DOBDO({\r6/t0/t2/s4/out_reg_n_16 ,\r6/t0/t2/s4/out_reg_n_17 ,\r6/t0/t2/s4/out_reg_n_18 ,\r6/t0/t2/s4/out_reg_n_19 ,\r6/t0/t2/s4/out_reg_n_20 ,\r6/t0/t2/s4/out_reg_n_21 ,\r6/t0/t2/s4/out_reg_n_22 ,\r6/t0/t2/s4/out_reg_n_23 ,\r6/t0/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r6/t1/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[95:88],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[87:80],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r6/t1/t0/s0/out_reg_n_0 ,\r6/t1/t0/s0/out_reg_n_1 ,\r6/t1/t0/s0/out_reg_n_2 ,\r6/t1/t0/s0/out_reg_n_3 ,\r6/t1/t0/s0/out_reg_n_4 ,\r6/t1/t0/s0/out_reg_n_5 ,\r6/t1/t0/s0/out_reg_n_6 ,\r6/t1/t0/s0/out_reg_n_7 ,\r6/t1/t0/p_0_in }),
        .DOBDO({\r6/t1/t0/s0/out_reg_n_16 ,\r6/t1/t0/s0/out_reg_n_17 ,\r6/t1/t0/s0/out_reg_n_18 ,\r6/t1/t0/s0/out_reg_n_19 ,\r6/t1/t0/s0/out_reg_n_20 ,\r6/t1/t0/s0/out_reg_n_21 ,\r6/t1/t0/s0/out_reg_n_22 ,\r6/t1/t0/s0/out_reg_n_23 ,\r6/t1/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r6/t1/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[95:88],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[87:80],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r6/t1/t0/s4/out_reg_n_0 ,\r6/t1/t0/s4/out_reg_n_1 ,\r6/t1/t0/s4/out_reg_n_2 ,\r6/t1/t0/s4/out_reg_n_3 ,\r6/t1/t0/s4/out_reg_n_4 ,\r6/t1/t0/s4/out_reg_n_5 ,\r6/t1/t0/s4/out_reg_n_6 ,\r6/t1/t0/s4/out_reg_n_7 ,\r6/t1/t0/p_1_in }),
        .DOBDO({\r6/t1/t0/s4/out_reg_n_16 ,\r6/t1/t0/s4/out_reg_n_17 ,\r6/t1/t0/s4/out_reg_n_18 ,\r6/t1/t0/s4/out_reg_n_19 ,\r6/t1/t0/s4/out_reg_n_20 ,\r6/t1/t0/s4/out_reg_n_21 ,\r6/t1/t0/s4/out_reg_n_22 ,\r6/t1/t0/s4/out_reg_n_23 ,\r6/t1/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r6/t1/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[79:72],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[71:64],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r6/t1/t2/s0/out_reg_n_0 ,\r6/t1/t2/s0/out_reg_n_1 ,\r6/t1/t2/s0/out_reg_n_2 ,\r6/t1/t2/s0/out_reg_n_3 ,\r6/t1/t2/s0/out_reg_n_4 ,\r6/t1/t2/s0/out_reg_n_5 ,\r6/t1/t2/s0/out_reg_n_6 ,\r6/t1/t2/s0/out_reg_n_7 ,\r6/t1/t2/p_0_in }),
        .DOBDO({\r6/t1/t2/s0/out_reg_n_16 ,\r6/t1/t2/s0/out_reg_n_17 ,\r6/t1/t2/s0/out_reg_n_18 ,\r6/t1/t2/s0/out_reg_n_19 ,\r6/t1/t2/s0/out_reg_n_20 ,\r6/t1/t2/s0/out_reg_n_21 ,\r6/t1/t2/s0/out_reg_n_22 ,\r6/t1/t2/s0/out_reg_n_23 ,\r6/t1/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r6/t1/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[79:72],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[71:64],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r6/t1/t2/s4/out_reg_n_0 ,\r6/t1/t2/s4/out_reg_n_1 ,\r6/t1/t2/s4/out_reg_n_2 ,\r6/t1/t2/s4/out_reg_n_3 ,\r6/t1/t2/s4/out_reg_n_4 ,\r6/t1/t2/s4/out_reg_n_5 ,\r6/t1/t2/s4/out_reg_n_6 ,\r6/t1/t2/s4/out_reg_n_7 ,\r6/t1/t2/p_1_in }),
        .DOBDO({\r6/t1/t2/s4/out_reg_n_16 ,\r6/t1/t2/s4/out_reg_n_17 ,\r6/t1/t2/s4/out_reg_n_18 ,\r6/t1/t2/s4/out_reg_n_19 ,\r6/t1/t2/s4/out_reg_n_20 ,\r6/t1/t2/s4/out_reg_n_21 ,\r6/t1/t2/s4/out_reg_n_22 ,\r6/t1/t2/s4/out_reg_n_23 ,\r6/t1/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r6/t2/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[63:56],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[55:48],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r6/t2/t0/s0/out_reg_n_0 ,\r6/t2/t0/s0/out_reg_n_1 ,\r6/t2/t0/s0/out_reg_n_2 ,\r6/t2/t0/s0/out_reg_n_3 ,\r6/t2/t0/s0/out_reg_n_4 ,\r6/t2/t0/s0/out_reg_n_5 ,\r6/t2/t0/s0/out_reg_n_6 ,\r6/t2/t0/s0/out_reg_n_7 ,\r6/t2/t0/p_0_in }),
        .DOBDO({\r6/t2/t0/s0/out_reg_n_16 ,\r6/t2/t0/s0/out_reg_n_17 ,\r6/t2/t0/s0/out_reg_n_18 ,\r6/t2/t0/s0/out_reg_n_19 ,\r6/t2/t0/s0/out_reg_n_20 ,\r6/t2/t0/s0/out_reg_n_21 ,\r6/t2/t0/s0/out_reg_n_22 ,\r6/t2/t0/s0/out_reg_n_23 ,\r6/t2/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r6/t2/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[63:56],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[55:48],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r6/t2/t0/s4/out_reg_n_0 ,\r6/t2/t0/s4/out_reg_n_1 ,\r6/t2/t0/s4/out_reg_n_2 ,\r6/t2/t0/s4/out_reg_n_3 ,\r6/t2/t0/s4/out_reg_n_4 ,\r6/t2/t0/s4/out_reg_n_5 ,\r6/t2/t0/s4/out_reg_n_6 ,\r6/t2/t0/s4/out_reg_n_7 ,\r6/t2/t0/p_1_in }),
        .DOBDO({\r6/t2/t0/s4/out_reg_n_16 ,\r6/t2/t0/s4/out_reg_n_17 ,\r6/t2/t0/s4/out_reg_n_18 ,\r6/t2/t0/s4/out_reg_n_19 ,\r6/t2/t0/s4/out_reg_n_20 ,\r6/t2/t0/s4/out_reg_n_21 ,\r6/t2/t0/s4/out_reg_n_22 ,\r6/t2/t0/s4/out_reg_n_23 ,\r6/t2/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r6/t2/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[47:40],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[39:32],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r6/t2/t2/s0/out_reg_n_0 ,\r6/t2/t2/s0/out_reg_n_1 ,\r6/t2/t2/s0/out_reg_n_2 ,\r6/t2/t2/s0/out_reg_n_3 ,\r6/t2/t2/s0/out_reg_n_4 ,\r6/t2/t2/s0/out_reg_n_5 ,\r6/t2/t2/s0/out_reg_n_6 ,\r6/t2/t2/s0/out_reg_n_7 ,\r6/t2/t2/p_0_in }),
        .DOBDO({\r6/t2/t2/s0/out_reg_n_16 ,\r6/t2/t2/s0/out_reg_n_17 ,\r6/t2/t2/s0/out_reg_n_18 ,\r6/t2/t2/s0/out_reg_n_19 ,\r6/t2/t2/s0/out_reg_n_20 ,\r6/t2/t2/s0/out_reg_n_21 ,\r6/t2/t2/s0/out_reg_n_22 ,\r6/t2/t2/s0/out_reg_n_23 ,\r6/t2/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r6/t2/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[47:40],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[39:32],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r6/t2/t2/s4/out_reg_n_0 ,\r6/t2/t2/s4/out_reg_n_1 ,\r6/t2/t2/s4/out_reg_n_2 ,\r6/t2/t2/s4/out_reg_n_3 ,\r6/t2/t2/s4/out_reg_n_4 ,\r6/t2/t2/s4/out_reg_n_5 ,\r6/t2/t2/s4/out_reg_n_6 ,\r6/t2/t2/s4/out_reg_n_7 ,\r6/t2/t2/p_1_in }),
        .DOBDO({\r6/t2/t2/s4/out_reg_n_16 ,\r6/t2/t2/s4/out_reg_n_17 ,\r6/t2/t2/s4/out_reg_n_18 ,\r6/t2/t2/s4/out_reg_n_19 ,\r6/t2/t2/s4/out_reg_n_20 ,\r6/t2/t2/s4/out_reg_n_21 ,\r6/t2/t2/s4/out_reg_n_22 ,\r6/t2/t2/s4/out_reg_n_23 ,\r6/t2/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r6/t3/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r6/t3/t0/s0/out_reg_n_0 ,\r6/t3/t0/s0/out_reg_n_1 ,\r6/t3/t0/s0/out_reg_n_2 ,\r6/t3/t0/s0/out_reg_n_3 ,\r6/t3/t0/s0/out_reg_n_4 ,\r6/t3/t0/s0/out_reg_n_5 ,\r6/t3/t0/s0/out_reg_n_6 ,\r6/t3/t0/s0/out_reg_n_7 ,\r6/t3/t0/p_0_in }),
        .DOBDO({\r6/t3/t0/s0/out_reg_n_16 ,\r6/t3/t0/s0/out_reg_n_17 ,\r6/t3/t0/s0/out_reg_n_18 ,\r6/t3/t0/s0/out_reg_n_19 ,\r6/t3/t0/s0/out_reg_n_20 ,\r6/t3/t0/s0/out_reg_n_21 ,\r6/t3/t0/s0/out_reg_n_22 ,\r6/t3/t0/s0/out_reg_n_23 ,\r6/t3/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r6/t3/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r6/t3/t0/s4/out_reg_n_0 ,\r6/t3/t0/s4/out_reg_n_1 ,\r6/t3/t0/s4/out_reg_n_2 ,\r6/t3/t0/s4/out_reg_n_3 ,\r6/t3/t0/s4/out_reg_n_4 ,\r6/t3/t0/s4/out_reg_n_5 ,\r6/t3/t0/s4/out_reg_n_6 ,\r6/t3/t0/s4/out_reg_n_7 ,\r6/t3/t0/p_1_in }),
        .DOBDO({\r6/t3/t0/s4/out_reg_n_16 ,\r6/t3/t0/s4/out_reg_n_17 ,\r6/t3/t0/s4/out_reg_n_18 ,\r6/t3/t0/s4/out_reg_n_19 ,\r6/t3/t0/s4/out_reg_n_20 ,\r6/t3/t0/s4/out_reg_n_21 ,\r6/t3/t0/s4/out_reg_n_22 ,\r6/t3/t0/s4/out_reg_n_23 ,\r6/t3/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r6/t3/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r6/t3/t2/s0/out_reg_n_0 ,\r6/t3/t2/s0/out_reg_n_1 ,\r6/t3/t2/s0/out_reg_n_2 ,\r6/t3/t2/s0/out_reg_n_3 ,\r6/t3/t2/s0/out_reg_n_4 ,\r6/t3/t2/s0/out_reg_n_5 ,\r6/t3/t2/s0/out_reg_n_6 ,\r6/t3/t2/s0/out_reg_n_7 ,\r6/t3/t2/p_0_in }),
        .DOBDO({\r6/t3/t2/s0/out_reg_n_16 ,\r6/t3/t2/s0/out_reg_n_17 ,\r6/t3/t2/s0/out_reg_n_18 ,\r6/t3/t2/s0/out_reg_n_19 ,\r6/t3/t2/s0/out_reg_n_20 ,\r6/t3/t2/s0/out_reg_n_21 ,\r6/t3/t2/s0/out_reg_n_22 ,\r6/t3/t2/s0/out_reg_n_23 ,\r6/t3/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r6/t3/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s5[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r6/t3/t2/s4/out_reg_n_0 ,\r6/t3/t2/s4/out_reg_n_1 ,\r6/t3/t2/s4/out_reg_n_2 ,\r6/t3/t2/s4/out_reg_n_3 ,\r6/t3/t2/s4/out_reg_n_4 ,\r6/t3/t2/s4/out_reg_n_5 ,\r6/t3/t2/s4/out_reg_n_6 ,\r6/t3/t2/s4/out_reg_n_7 ,\r6/t3/t2/p_1_in }),
        .DOBDO({\r6/t3/t2/s4/out_reg_n_16 ,\r6/t3/t2/s4/out_reg_n_17 ,\r6/t3/t2/s4/out_reg_n_18 ,\r6/t3/t2/s4/out_reg_n_19 ,\r6/t3/t2/s4/out_reg_n_20 ,\r6/t3/t2/s4/out_reg_n_21 ,\r6/t3/t2/s4/out_reg_n_22 ,\r6/t3/t2/s4/out_reg_n_23 ,\r6/t3/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [0]),
        .Q(s7[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[100] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [100]),
        .Q(s7[100]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[101] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [101]),
        .Q(s7[101]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[102] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [102]),
        .Q(s7[102]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[103] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [103]),
        .Q(s7[103]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[104] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [104]),
        .Q(s7[104]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[105] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [105]),
        .Q(s7[105]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[106] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [106]),
        .Q(s7[106]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[107] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [107]),
        .Q(s7[107]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[108] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [108]),
        .Q(s7[108]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[109] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [109]),
        .Q(s7[109]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [10]),
        .Q(s7[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[110] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [110]),
        .Q(s7[110]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[111] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [111]),
        .Q(s7[111]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[112] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [112]),
        .Q(s7[112]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[113] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [113]),
        .Q(s7[113]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[114] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [114]),
        .Q(s7[114]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[115] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [115]),
        .Q(s7[115]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[116] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [116]),
        .Q(s7[116]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[117] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [117]),
        .Q(s7[117]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[118] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [118]),
        .Q(s7[118]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[119] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [119]),
        .Q(s7[119]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [11]),
        .Q(s7[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[120] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [120]),
        .Q(s7[120]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[121] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [121]),
        .Q(s7[121]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[122] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [122]),
        .Q(s7[122]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[123] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [123]),
        .Q(s7[123]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[124] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [124]),
        .Q(s7[124]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[125] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [125]),
        .Q(s7[125]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[126] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [126]),
        .Q(s7[126]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[127] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [127]),
        .Q(s7[127]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [12]),
        .Q(s7[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [13]),
        .Q(s7[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [14]),
        .Q(s7[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [15]),
        .Q(s7[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [16]),
        .Q(s7[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [17]),
        .Q(s7[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [18]),
        .Q(s7[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [19]),
        .Q(s7[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [1]),
        .Q(s7[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [20]),
        .Q(s7[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [21]),
        .Q(s7[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [22]),
        .Q(s7[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [23]),
        .Q(s7[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [24]),
        .Q(s7[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [25]),
        .Q(s7[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [26]),
        .Q(s7[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [27]),
        .Q(s7[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [28]),
        .Q(s7[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [29]),
        .Q(s7[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [2]),
        .Q(s7[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [30]),
        .Q(s7[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [31]),
        .Q(s7[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [32]),
        .Q(s7[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [33]),
        .Q(s7[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [34]),
        .Q(s7[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [35]),
        .Q(s7[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [36]),
        .Q(s7[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [37]),
        .Q(s7[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [38]),
        .Q(s7[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [39]),
        .Q(s7[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [3]),
        .Q(s7[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [40]),
        .Q(s7[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [41]),
        .Q(s7[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [42]),
        .Q(s7[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [43]),
        .Q(s7[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [44]),
        .Q(s7[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [45]),
        .Q(s7[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [46]),
        .Q(s7[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [47]),
        .Q(s7[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [48]),
        .Q(s7[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [49]),
        .Q(s7[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [4]),
        .Q(s7[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [50]),
        .Q(s7[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [51]),
        .Q(s7[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [52]),
        .Q(s7[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [53]),
        .Q(s7[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [54]),
        .Q(s7[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [55]),
        .Q(s7[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [56]),
        .Q(s7[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [57]),
        .Q(s7[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [58]),
        .Q(s7[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [59]),
        .Q(s7[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [5]),
        .Q(s7[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [60]),
        .Q(s7[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [61]),
        .Q(s7[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [62]),
        .Q(s7[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [63]),
        .Q(s7[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[64] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [64]),
        .Q(s7[64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[65] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [65]),
        .Q(s7[65]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[66] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [66]),
        .Q(s7[66]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[67] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [67]),
        .Q(s7[67]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[68] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [68]),
        .Q(s7[68]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[69] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [69]),
        .Q(s7[69]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [6]),
        .Q(s7[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[70] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [70]),
        .Q(s7[70]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[71] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [71]),
        .Q(s7[71]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[72] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [72]),
        .Q(s7[72]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[73] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [73]),
        .Q(s7[73]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[74] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [74]),
        .Q(s7[74]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[75] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [75]),
        .Q(s7[75]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[76] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [76]),
        .Q(s7[76]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[77] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [77]),
        .Q(s7[77]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[78] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [78]),
        .Q(s7[78]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[79] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [79]),
        .Q(s7[79]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [7]),
        .Q(s7[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[80] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [80]),
        .Q(s7[80]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[81] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [81]),
        .Q(s7[81]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[82] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [82]),
        .Q(s7[82]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[83] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [83]),
        .Q(s7[83]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[84] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [84]),
        .Q(s7[84]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[85] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [85]),
        .Q(s7[85]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[86] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [86]),
        .Q(s7[86]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[87] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [87]),
        .Q(s7[87]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[88] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [88]),
        .Q(s7[88]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[89] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [89]),
        .Q(s7[89]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [8]),
        .Q(s7[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[90] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [90]),
        .Q(s7[90]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[91] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [91]),
        .Q(s7[91]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[92] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [92]),
        .Q(s7[92]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[93] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [93]),
        .Q(s7[93]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[94] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [94]),
        .Q(s7[94]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[95] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [95]),
        .Q(s7[95]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[96] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [96]),
        .Q(s7[96]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[97] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [97]),
        .Q(s7[97]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[98] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [98]),
        .Q(s7[98]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[99] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [99]),
        .Q(s7[99]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r7/state_out_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r7/p_0_out [9]),
        .Q(s7[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r7/t0/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[127:120],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[119:112],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r7/t0/t0/s0/out_reg_n_0 ,\r7/t0/t0/s0/out_reg_n_1 ,\r7/t0/t0/s0/out_reg_n_2 ,\r7/t0/t0/s0/out_reg_n_3 ,\r7/t0/t0/s0/out_reg_n_4 ,\r7/t0/t0/s0/out_reg_n_5 ,\r7/t0/t0/s0/out_reg_n_6 ,\r7/t0/t0/s0/out_reg_n_7 ,\r7/t0/t0/p_0_in }),
        .DOBDO({\r7/t0/t0/s0/out_reg_n_16 ,\r7/t0/t0/s0/out_reg_n_17 ,\r7/t0/t0/s0/out_reg_n_18 ,\r7/t0/t0/s0/out_reg_n_19 ,\r7/t0/t0/s0/out_reg_n_20 ,\r7/t0/t0/s0/out_reg_n_21 ,\r7/t0/t0/s0/out_reg_n_22 ,\r7/t0/t0/s0/out_reg_n_23 ,\r7/t0/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r7/t0/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[127:120],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[119:112],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r7/t0/t0/s4/out_reg_n_0 ,\r7/t0/t0/s4/out_reg_n_1 ,\r7/t0/t0/s4/out_reg_n_2 ,\r7/t0/t0/s4/out_reg_n_3 ,\r7/t0/t0/s4/out_reg_n_4 ,\r7/t0/t0/s4/out_reg_n_5 ,\r7/t0/t0/s4/out_reg_n_6 ,\r7/t0/t0/s4/out_reg_n_7 ,\r7/t0/t0/p_1_in }),
        .DOBDO({\r7/t0/t0/s4/out_reg_n_16 ,\r7/t0/t0/s4/out_reg_n_17 ,\r7/t0/t0/s4/out_reg_n_18 ,\r7/t0/t0/s4/out_reg_n_19 ,\r7/t0/t0/s4/out_reg_n_20 ,\r7/t0/t0/s4/out_reg_n_21 ,\r7/t0/t0/s4/out_reg_n_22 ,\r7/t0/t0/s4/out_reg_n_23 ,\r7/t0/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r7/t0/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[111:104],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[103:96],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r7/t0/t2/s0/out_reg_n_0 ,\r7/t0/t2/s0/out_reg_n_1 ,\r7/t0/t2/s0/out_reg_n_2 ,\r7/t0/t2/s0/out_reg_n_3 ,\r7/t0/t2/s0/out_reg_n_4 ,\r7/t0/t2/s0/out_reg_n_5 ,\r7/t0/t2/s0/out_reg_n_6 ,\r7/t0/t2/s0/out_reg_n_7 ,\r7/t0/t2/p_0_in }),
        .DOBDO({\r7/t0/t2/s0/out_reg_n_16 ,\r7/t0/t2/s0/out_reg_n_17 ,\r7/t0/t2/s0/out_reg_n_18 ,\r7/t0/t2/s0/out_reg_n_19 ,\r7/t0/t2/s0/out_reg_n_20 ,\r7/t0/t2/s0/out_reg_n_21 ,\r7/t0/t2/s0/out_reg_n_22 ,\r7/t0/t2/s0/out_reg_n_23 ,\r7/t0/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r7/t0/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[111:104],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[103:96],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r7/t0/t2/s4/out_reg_n_0 ,\r7/t0/t2/s4/out_reg_n_1 ,\r7/t0/t2/s4/out_reg_n_2 ,\r7/t0/t2/s4/out_reg_n_3 ,\r7/t0/t2/s4/out_reg_n_4 ,\r7/t0/t2/s4/out_reg_n_5 ,\r7/t0/t2/s4/out_reg_n_6 ,\r7/t0/t2/s4/out_reg_n_7 ,\r7/t0/t2/p_1_in }),
        .DOBDO({\r7/t0/t2/s4/out_reg_n_16 ,\r7/t0/t2/s4/out_reg_n_17 ,\r7/t0/t2/s4/out_reg_n_18 ,\r7/t0/t2/s4/out_reg_n_19 ,\r7/t0/t2/s4/out_reg_n_20 ,\r7/t0/t2/s4/out_reg_n_21 ,\r7/t0/t2/s4/out_reg_n_22 ,\r7/t0/t2/s4/out_reg_n_23 ,\r7/t0/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r7/t1/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[95:88],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[87:80],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r7/t1/t0/s0/out_reg_n_0 ,\r7/t1/t0/s0/out_reg_n_1 ,\r7/t1/t0/s0/out_reg_n_2 ,\r7/t1/t0/s0/out_reg_n_3 ,\r7/t1/t0/s0/out_reg_n_4 ,\r7/t1/t0/s0/out_reg_n_5 ,\r7/t1/t0/s0/out_reg_n_6 ,\r7/t1/t0/s0/out_reg_n_7 ,\r7/t1/t0/p_0_in }),
        .DOBDO({\r7/t1/t0/s0/out_reg_n_16 ,\r7/t1/t0/s0/out_reg_n_17 ,\r7/t1/t0/s0/out_reg_n_18 ,\r7/t1/t0/s0/out_reg_n_19 ,\r7/t1/t0/s0/out_reg_n_20 ,\r7/t1/t0/s0/out_reg_n_21 ,\r7/t1/t0/s0/out_reg_n_22 ,\r7/t1/t0/s0/out_reg_n_23 ,\r7/t1/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r7/t1/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[95:88],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[87:80],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r7/t1/t0/s4/out_reg_n_0 ,\r7/t1/t0/s4/out_reg_n_1 ,\r7/t1/t0/s4/out_reg_n_2 ,\r7/t1/t0/s4/out_reg_n_3 ,\r7/t1/t0/s4/out_reg_n_4 ,\r7/t1/t0/s4/out_reg_n_5 ,\r7/t1/t0/s4/out_reg_n_6 ,\r7/t1/t0/s4/out_reg_n_7 ,\r7/t1/t0/p_1_in }),
        .DOBDO({\r7/t1/t0/s4/out_reg_n_16 ,\r7/t1/t0/s4/out_reg_n_17 ,\r7/t1/t0/s4/out_reg_n_18 ,\r7/t1/t0/s4/out_reg_n_19 ,\r7/t1/t0/s4/out_reg_n_20 ,\r7/t1/t0/s4/out_reg_n_21 ,\r7/t1/t0/s4/out_reg_n_22 ,\r7/t1/t0/s4/out_reg_n_23 ,\r7/t1/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r7/t1/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[79:72],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[71:64],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r7/t1/t2/s0/out_reg_n_0 ,\r7/t1/t2/s0/out_reg_n_1 ,\r7/t1/t2/s0/out_reg_n_2 ,\r7/t1/t2/s0/out_reg_n_3 ,\r7/t1/t2/s0/out_reg_n_4 ,\r7/t1/t2/s0/out_reg_n_5 ,\r7/t1/t2/s0/out_reg_n_6 ,\r7/t1/t2/s0/out_reg_n_7 ,\r7/t1/t2/p_0_in }),
        .DOBDO({\r7/t1/t2/s0/out_reg_n_16 ,\r7/t1/t2/s0/out_reg_n_17 ,\r7/t1/t2/s0/out_reg_n_18 ,\r7/t1/t2/s0/out_reg_n_19 ,\r7/t1/t2/s0/out_reg_n_20 ,\r7/t1/t2/s0/out_reg_n_21 ,\r7/t1/t2/s0/out_reg_n_22 ,\r7/t1/t2/s0/out_reg_n_23 ,\r7/t1/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r7/t1/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[79:72],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[71:64],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r7/t1/t2/s4/out_reg_n_0 ,\r7/t1/t2/s4/out_reg_n_1 ,\r7/t1/t2/s4/out_reg_n_2 ,\r7/t1/t2/s4/out_reg_n_3 ,\r7/t1/t2/s4/out_reg_n_4 ,\r7/t1/t2/s4/out_reg_n_5 ,\r7/t1/t2/s4/out_reg_n_6 ,\r7/t1/t2/s4/out_reg_n_7 ,\r7/t1/t2/p_1_in }),
        .DOBDO({\r7/t1/t2/s4/out_reg_n_16 ,\r7/t1/t2/s4/out_reg_n_17 ,\r7/t1/t2/s4/out_reg_n_18 ,\r7/t1/t2/s4/out_reg_n_19 ,\r7/t1/t2/s4/out_reg_n_20 ,\r7/t1/t2/s4/out_reg_n_21 ,\r7/t1/t2/s4/out_reg_n_22 ,\r7/t1/t2/s4/out_reg_n_23 ,\r7/t1/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r7/t2/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[63:56],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[55:48],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r7/t2/t0/s0/out_reg_n_0 ,\r7/t2/t0/s0/out_reg_n_1 ,\r7/t2/t0/s0/out_reg_n_2 ,\r7/t2/t0/s0/out_reg_n_3 ,\r7/t2/t0/s0/out_reg_n_4 ,\r7/t2/t0/s0/out_reg_n_5 ,\r7/t2/t0/s0/out_reg_n_6 ,\r7/t2/t0/s0/out_reg_n_7 ,\r7/t2/t0/p_0_in }),
        .DOBDO({\r7/t2/t0/s0/out_reg_n_16 ,\r7/t2/t0/s0/out_reg_n_17 ,\r7/t2/t0/s0/out_reg_n_18 ,\r7/t2/t0/s0/out_reg_n_19 ,\r7/t2/t0/s0/out_reg_n_20 ,\r7/t2/t0/s0/out_reg_n_21 ,\r7/t2/t0/s0/out_reg_n_22 ,\r7/t2/t0/s0/out_reg_n_23 ,\r7/t2/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r7/t2/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[63:56],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[55:48],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r7/t2/t0/s4/out_reg_n_0 ,\r7/t2/t0/s4/out_reg_n_1 ,\r7/t2/t0/s4/out_reg_n_2 ,\r7/t2/t0/s4/out_reg_n_3 ,\r7/t2/t0/s4/out_reg_n_4 ,\r7/t2/t0/s4/out_reg_n_5 ,\r7/t2/t0/s4/out_reg_n_6 ,\r7/t2/t0/s4/out_reg_n_7 ,\r7/t2/t0/p_1_in }),
        .DOBDO({\r7/t2/t0/s4/out_reg_n_16 ,\r7/t2/t0/s4/out_reg_n_17 ,\r7/t2/t0/s4/out_reg_n_18 ,\r7/t2/t0/s4/out_reg_n_19 ,\r7/t2/t0/s4/out_reg_n_20 ,\r7/t2/t0/s4/out_reg_n_21 ,\r7/t2/t0/s4/out_reg_n_22 ,\r7/t2/t0/s4/out_reg_n_23 ,\r7/t2/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r7/t2/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[47:40],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[39:32],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r7/t2/t2/s0/out_reg_n_0 ,\r7/t2/t2/s0/out_reg_n_1 ,\r7/t2/t2/s0/out_reg_n_2 ,\r7/t2/t2/s0/out_reg_n_3 ,\r7/t2/t2/s0/out_reg_n_4 ,\r7/t2/t2/s0/out_reg_n_5 ,\r7/t2/t2/s0/out_reg_n_6 ,\r7/t2/t2/s0/out_reg_n_7 ,\r7/t2/t2/p_0_in }),
        .DOBDO({\r7/t2/t2/s0/out_reg_n_16 ,\r7/t2/t2/s0/out_reg_n_17 ,\r7/t2/t2/s0/out_reg_n_18 ,\r7/t2/t2/s0/out_reg_n_19 ,\r7/t2/t2/s0/out_reg_n_20 ,\r7/t2/t2/s0/out_reg_n_21 ,\r7/t2/t2/s0/out_reg_n_22 ,\r7/t2/t2/s0/out_reg_n_23 ,\r7/t2/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r7/t2/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[47:40],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[39:32],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r7/t2/t2/s4/out_reg_n_0 ,\r7/t2/t2/s4/out_reg_n_1 ,\r7/t2/t2/s4/out_reg_n_2 ,\r7/t2/t2/s4/out_reg_n_3 ,\r7/t2/t2/s4/out_reg_n_4 ,\r7/t2/t2/s4/out_reg_n_5 ,\r7/t2/t2/s4/out_reg_n_6 ,\r7/t2/t2/s4/out_reg_n_7 ,\r7/t2/t2/p_1_in }),
        .DOBDO({\r7/t2/t2/s4/out_reg_n_16 ,\r7/t2/t2/s4/out_reg_n_17 ,\r7/t2/t2/s4/out_reg_n_18 ,\r7/t2/t2/s4/out_reg_n_19 ,\r7/t2/t2/s4/out_reg_n_20 ,\r7/t2/t2/s4/out_reg_n_21 ,\r7/t2/t2/s4/out_reg_n_22 ,\r7/t2/t2/s4/out_reg_n_23 ,\r7/t2/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r7/t3/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r7/t3/t0/s0/out_reg_n_0 ,\r7/t3/t0/s0/out_reg_n_1 ,\r7/t3/t0/s0/out_reg_n_2 ,\r7/t3/t0/s0/out_reg_n_3 ,\r7/t3/t0/s0/out_reg_n_4 ,\r7/t3/t0/s0/out_reg_n_5 ,\r7/t3/t0/s0/out_reg_n_6 ,\r7/t3/t0/s0/out_reg_n_7 ,\r7/t3/t0/p_0_in }),
        .DOBDO({\r7/t3/t0/s0/out_reg_n_16 ,\r7/t3/t0/s0/out_reg_n_17 ,\r7/t3/t0/s0/out_reg_n_18 ,\r7/t3/t0/s0/out_reg_n_19 ,\r7/t3/t0/s0/out_reg_n_20 ,\r7/t3/t0/s0/out_reg_n_21 ,\r7/t3/t0/s0/out_reg_n_22 ,\r7/t3/t0/s0/out_reg_n_23 ,\r7/t3/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r7/t3/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r7/t3/t0/s4/out_reg_n_0 ,\r7/t3/t0/s4/out_reg_n_1 ,\r7/t3/t0/s4/out_reg_n_2 ,\r7/t3/t0/s4/out_reg_n_3 ,\r7/t3/t0/s4/out_reg_n_4 ,\r7/t3/t0/s4/out_reg_n_5 ,\r7/t3/t0/s4/out_reg_n_6 ,\r7/t3/t0/s4/out_reg_n_7 ,\r7/t3/t0/p_1_in }),
        .DOBDO({\r7/t3/t0/s4/out_reg_n_16 ,\r7/t3/t0/s4/out_reg_n_17 ,\r7/t3/t0/s4/out_reg_n_18 ,\r7/t3/t0/s4/out_reg_n_19 ,\r7/t3/t0/s4/out_reg_n_20 ,\r7/t3/t0/s4/out_reg_n_21 ,\r7/t3/t0/s4/out_reg_n_22 ,\r7/t3/t0/s4/out_reg_n_23 ,\r7/t3/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r7/t3/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r7/t3/t2/s0/out_reg_n_0 ,\r7/t3/t2/s0/out_reg_n_1 ,\r7/t3/t2/s0/out_reg_n_2 ,\r7/t3/t2/s0/out_reg_n_3 ,\r7/t3/t2/s0/out_reg_n_4 ,\r7/t3/t2/s0/out_reg_n_5 ,\r7/t3/t2/s0/out_reg_n_6 ,\r7/t3/t2/s0/out_reg_n_7 ,\r7/t3/t2/p_0_in }),
        .DOBDO({\r7/t3/t2/s0/out_reg_n_16 ,\r7/t3/t2/s0/out_reg_n_17 ,\r7/t3/t2/s0/out_reg_n_18 ,\r7/t3/t2/s0/out_reg_n_19 ,\r7/t3/t2/s0/out_reg_n_20 ,\r7/t3/t2/s0/out_reg_n_21 ,\r7/t3/t2/s0/out_reg_n_22 ,\r7/t3/t2/s0/out_reg_n_23 ,\r7/t3/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r7/t3/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s6[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r7/t3/t2/s4/out_reg_n_0 ,\r7/t3/t2/s4/out_reg_n_1 ,\r7/t3/t2/s4/out_reg_n_2 ,\r7/t3/t2/s4/out_reg_n_3 ,\r7/t3/t2/s4/out_reg_n_4 ,\r7/t3/t2/s4/out_reg_n_5 ,\r7/t3/t2/s4/out_reg_n_6 ,\r7/t3/t2/s4/out_reg_n_7 ,\r7/t3/t2/p_1_in }),
        .DOBDO({\r7/t3/t2/s4/out_reg_n_16 ,\r7/t3/t2/s4/out_reg_n_17 ,\r7/t3/t2/s4/out_reg_n_18 ,\r7/t3/t2/s4/out_reg_n_19 ,\r7/t3/t2/s4/out_reg_n_20 ,\r7/t3/t2/s4/out_reg_n_21 ,\r7/t3/t2/s4/out_reg_n_22 ,\r7/t3/t2/s4/out_reg_n_23 ,\r7/t3/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [0]),
        .Q(s8[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[100] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [100]),
        .Q(s8[100]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[101] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [101]),
        .Q(s8[101]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[102] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [102]),
        .Q(s8[102]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[103] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [103]),
        .Q(s8[103]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[104] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [104]),
        .Q(s8[104]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[105] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [105]),
        .Q(s8[105]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[106] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [106]),
        .Q(s8[106]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[107] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [107]),
        .Q(s8[107]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[108] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [108]),
        .Q(s8[108]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[109] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [109]),
        .Q(s8[109]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [10]),
        .Q(s8[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[110] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [110]),
        .Q(s8[110]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[111] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [111]),
        .Q(s8[111]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[112] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [112]),
        .Q(s8[112]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[113] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [113]),
        .Q(s8[113]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[114] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [114]),
        .Q(s8[114]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[115] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [115]),
        .Q(s8[115]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[116] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [116]),
        .Q(s8[116]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[117] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [117]),
        .Q(s8[117]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[118] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [118]),
        .Q(s8[118]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[119] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [119]),
        .Q(s8[119]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [11]),
        .Q(s8[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[120] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [120]),
        .Q(s8[120]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[121] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [121]),
        .Q(s8[121]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[122] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [122]),
        .Q(s8[122]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[123] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [123]),
        .Q(s8[123]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[124] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [124]),
        .Q(s8[124]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[125] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [125]),
        .Q(s8[125]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[126] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [126]),
        .Q(s8[126]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[127] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [127]),
        .Q(s8[127]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [12]),
        .Q(s8[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [13]),
        .Q(s8[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [14]),
        .Q(s8[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [15]),
        .Q(s8[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [16]),
        .Q(s8[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [17]),
        .Q(s8[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [18]),
        .Q(s8[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [19]),
        .Q(s8[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [1]),
        .Q(s8[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [20]),
        .Q(s8[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [21]),
        .Q(s8[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [22]),
        .Q(s8[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [23]),
        .Q(s8[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [24]),
        .Q(s8[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [25]),
        .Q(s8[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [26]),
        .Q(s8[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [27]),
        .Q(s8[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [28]),
        .Q(s8[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [29]),
        .Q(s8[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [2]),
        .Q(s8[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [30]),
        .Q(s8[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [31]),
        .Q(s8[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [32]),
        .Q(s8[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [33]),
        .Q(s8[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [34]),
        .Q(s8[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [35]),
        .Q(s8[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [36]),
        .Q(s8[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [37]),
        .Q(s8[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [38]),
        .Q(s8[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [39]),
        .Q(s8[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [3]),
        .Q(s8[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [40]),
        .Q(s8[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [41]),
        .Q(s8[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [42]),
        .Q(s8[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [43]),
        .Q(s8[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [44]),
        .Q(s8[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [45]),
        .Q(s8[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [46]),
        .Q(s8[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [47]),
        .Q(s8[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [48]),
        .Q(s8[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [49]),
        .Q(s8[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [4]),
        .Q(s8[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [50]),
        .Q(s8[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [51]),
        .Q(s8[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [52]),
        .Q(s8[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [53]),
        .Q(s8[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [54]),
        .Q(s8[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [55]),
        .Q(s8[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [56]),
        .Q(s8[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [57]),
        .Q(s8[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [58]),
        .Q(s8[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [59]),
        .Q(s8[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [5]),
        .Q(s8[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [60]),
        .Q(s8[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [61]),
        .Q(s8[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [62]),
        .Q(s8[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [63]),
        .Q(s8[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[64] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [64]),
        .Q(s8[64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[65] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [65]),
        .Q(s8[65]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[66] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [66]),
        .Q(s8[66]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[67] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [67]),
        .Q(s8[67]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[68] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [68]),
        .Q(s8[68]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[69] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [69]),
        .Q(s8[69]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [6]),
        .Q(s8[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[70] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [70]),
        .Q(s8[70]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[71] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [71]),
        .Q(s8[71]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[72] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [72]),
        .Q(s8[72]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[73] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [73]),
        .Q(s8[73]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[74] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [74]),
        .Q(s8[74]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[75] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [75]),
        .Q(s8[75]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[76] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [76]),
        .Q(s8[76]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[77] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [77]),
        .Q(s8[77]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[78] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [78]),
        .Q(s8[78]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[79] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [79]),
        .Q(s8[79]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [7]),
        .Q(s8[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[80] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [80]),
        .Q(s8[80]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[81] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [81]),
        .Q(s8[81]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[82] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [82]),
        .Q(s8[82]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[83] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [83]),
        .Q(s8[83]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[84] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [84]),
        .Q(s8[84]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[85] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [85]),
        .Q(s8[85]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[86] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [86]),
        .Q(s8[86]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[87] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [87]),
        .Q(s8[87]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[88] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [88]),
        .Q(s8[88]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[89] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [89]),
        .Q(s8[89]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [8]),
        .Q(s8[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[90] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [90]),
        .Q(s8[90]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[91] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [91]),
        .Q(s8[91]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[92] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [92]),
        .Q(s8[92]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[93] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [93]),
        .Q(s8[93]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[94] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [94]),
        .Q(s8[94]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[95] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [95]),
        .Q(s8[95]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[96] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [96]),
        .Q(s8[96]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[97] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [97]),
        .Q(s8[97]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[98] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [98]),
        .Q(s8[98]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[99] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [99]),
        .Q(s8[99]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r8/state_out_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r8/p_0_out [9]),
        .Q(s8[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r8/t0/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[127:120],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[119:112],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r8/t0/t0/s0/out_reg_n_0 ,\r8/t0/t0/s0/out_reg_n_1 ,\r8/t0/t0/s0/out_reg_n_2 ,\r8/t0/t0/s0/out_reg_n_3 ,\r8/t0/t0/s0/out_reg_n_4 ,\r8/t0/t0/s0/out_reg_n_5 ,\r8/t0/t0/s0/out_reg_n_6 ,\r8/t0/t0/s0/out_reg_n_7 ,\r8/t0/t0/p_0_in }),
        .DOBDO({\r8/t0/t0/s0/out_reg_n_16 ,\r8/t0/t0/s0/out_reg_n_17 ,\r8/t0/t0/s0/out_reg_n_18 ,\r8/t0/t0/s0/out_reg_n_19 ,\r8/t0/t0/s0/out_reg_n_20 ,\r8/t0/t0/s0/out_reg_n_21 ,\r8/t0/t0/s0/out_reg_n_22 ,\r8/t0/t0/s0/out_reg_n_23 ,\r8/t0/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r8/t0/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[127:120],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[119:112],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r8/t0/t0/s4/out_reg_n_0 ,\r8/t0/t0/s4/out_reg_n_1 ,\r8/t0/t0/s4/out_reg_n_2 ,\r8/t0/t0/s4/out_reg_n_3 ,\r8/t0/t0/s4/out_reg_n_4 ,\r8/t0/t0/s4/out_reg_n_5 ,\r8/t0/t0/s4/out_reg_n_6 ,\r8/t0/t0/s4/out_reg_n_7 ,\r8/t0/t0/p_1_in }),
        .DOBDO({\r8/t0/t0/s4/out_reg_n_16 ,\r8/t0/t0/s4/out_reg_n_17 ,\r8/t0/t0/s4/out_reg_n_18 ,\r8/t0/t0/s4/out_reg_n_19 ,\r8/t0/t0/s4/out_reg_n_20 ,\r8/t0/t0/s4/out_reg_n_21 ,\r8/t0/t0/s4/out_reg_n_22 ,\r8/t0/t0/s4/out_reg_n_23 ,\r8/t0/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r8/t0/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[111:104],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[103:96],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r8/t0/t2/s0/out_reg_n_0 ,\r8/t0/t2/s0/out_reg_n_1 ,\r8/t0/t2/s0/out_reg_n_2 ,\r8/t0/t2/s0/out_reg_n_3 ,\r8/t0/t2/s0/out_reg_n_4 ,\r8/t0/t2/s0/out_reg_n_5 ,\r8/t0/t2/s0/out_reg_n_6 ,\r8/t0/t2/s0/out_reg_n_7 ,\r8/t0/t2/p_0_in }),
        .DOBDO({\r8/t0/t2/s0/out_reg_n_16 ,\r8/t0/t2/s0/out_reg_n_17 ,\r8/t0/t2/s0/out_reg_n_18 ,\r8/t0/t2/s0/out_reg_n_19 ,\r8/t0/t2/s0/out_reg_n_20 ,\r8/t0/t2/s0/out_reg_n_21 ,\r8/t0/t2/s0/out_reg_n_22 ,\r8/t0/t2/s0/out_reg_n_23 ,\r8/t0/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r8/t0/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[111:104],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[103:96],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r8/t0/t2/s4/out_reg_n_0 ,\r8/t0/t2/s4/out_reg_n_1 ,\r8/t0/t2/s4/out_reg_n_2 ,\r8/t0/t2/s4/out_reg_n_3 ,\r8/t0/t2/s4/out_reg_n_4 ,\r8/t0/t2/s4/out_reg_n_5 ,\r8/t0/t2/s4/out_reg_n_6 ,\r8/t0/t2/s4/out_reg_n_7 ,\r8/t0/t2/p_1_in }),
        .DOBDO({\r8/t0/t2/s4/out_reg_n_16 ,\r8/t0/t2/s4/out_reg_n_17 ,\r8/t0/t2/s4/out_reg_n_18 ,\r8/t0/t2/s4/out_reg_n_19 ,\r8/t0/t2/s4/out_reg_n_20 ,\r8/t0/t2/s4/out_reg_n_21 ,\r8/t0/t2/s4/out_reg_n_22 ,\r8/t0/t2/s4/out_reg_n_23 ,\r8/t0/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r8/t1/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[95:88],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[87:80],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r8/t1/t0/s0/out_reg_n_0 ,\r8/t1/t0/s0/out_reg_n_1 ,\r8/t1/t0/s0/out_reg_n_2 ,\r8/t1/t0/s0/out_reg_n_3 ,\r8/t1/t0/s0/out_reg_n_4 ,\r8/t1/t0/s0/out_reg_n_5 ,\r8/t1/t0/s0/out_reg_n_6 ,\r8/t1/t0/s0/out_reg_n_7 ,\r8/t1/t0/p_0_in }),
        .DOBDO({\r8/t1/t0/s0/out_reg_n_16 ,\r8/t1/t0/s0/out_reg_n_17 ,\r8/t1/t0/s0/out_reg_n_18 ,\r8/t1/t0/s0/out_reg_n_19 ,\r8/t1/t0/s0/out_reg_n_20 ,\r8/t1/t0/s0/out_reg_n_21 ,\r8/t1/t0/s0/out_reg_n_22 ,\r8/t1/t0/s0/out_reg_n_23 ,\r8/t1/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r8/t1/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[95:88],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[87:80],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r8/t1/t0/s4/out_reg_n_0 ,\r8/t1/t0/s4/out_reg_n_1 ,\r8/t1/t0/s4/out_reg_n_2 ,\r8/t1/t0/s4/out_reg_n_3 ,\r8/t1/t0/s4/out_reg_n_4 ,\r8/t1/t0/s4/out_reg_n_5 ,\r8/t1/t0/s4/out_reg_n_6 ,\r8/t1/t0/s4/out_reg_n_7 ,\r8/t1/t0/p_1_in }),
        .DOBDO({\r8/t1/t0/s4/out_reg_n_16 ,\r8/t1/t0/s4/out_reg_n_17 ,\r8/t1/t0/s4/out_reg_n_18 ,\r8/t1/t0/s4/out_reg_n_19 ,\r8/t1/t0/s4/out_reg_n_20 ,\r8/t1/t0/s4/out_reg_n_21 ,\r8/t1/t0/s4/out_reg_n_22 ,\r8/t1/t0/s4/out_reg_n_23 ,\r8/t1/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r8/t1/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[79:72],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[71:64],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r8/t1/t2/s0/out_reg_n_0 ,\r8/t1/t2/s0/out_reg_n_1 ,\r8/t1/t2/s0/out_reg_n_2 ,\r8/t1/t2/s0/out_reg_n_3 ,\r8/t1/t2/s0/out_reg_n_4 ,\r8/t1/t2/s0/out_reg_n_5 ,\r8/t1/t2/s0/out_reg_n_6 ,\r8/t1/t2/s0/out_reg_n_7 ,\r8/t1/t2/p_0_in }),
        .DOBDO({\r8/t1/t2/s0/out_reg_n_16 ,\r8/t1/t2/s0/out_reg_n_17 ,\r8/t1/t2/s0/out_reg_n_18 ,\r8/t1/t2/s0/out_reg_n_19 ,\r8/t1/t2/s0/out_reg_n_20 ,\r8/t1/t2/s0/out_reg_n_21 ,\r8/t1/t2/s0/out_reg_n_22 ,\r8/t1/t2/s0/out_reg_n_23 ,\r8/t1/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r8/t1/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[79:72],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[71:64],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r8/t1/t2/s4/out_reg_n_0 ,\r8/t1/t2/s4/out_reg_n_1 ,\r8/t1/t2/s4/out_reg_n_2 ,\r8/t1/t2/s4/out_reg_n_3 ,\r8/t1/t2/s4/out_reg_n_4 ,\r8/t1/t2/s4/out_reg_n_5 ,\r8/t1/t2/s4/out_reg_n_6 ,\r8/t1/t2/s4/out_reg_n_7 ,\r8/t1/t2/p_1_in }),
        .DOBDO({\r8/t1/t2/s4/out_reg_n_16 ,\r8/t1/t2/s4/out_reg_n_17 ,\r8/t1/t2/s4/out_reg_n_18 ,\r8/t1/t2/s4/out_reg_n_19 ,\r8/t1/t2/s4/out_reg_n_20 ,\r8/t1/t2/s4/out_reg_n_21 ,\r8/t1/t2/s4/out_reg_n_22 ,\r8/t1/t2/s4/out_reg_n_23 ,\r8/t1/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r8/t2/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[63:56],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[55:48],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r8/t2/t0/s0/out_reg_n_0 ,\r8/t2/t0/s0/out_reg_n_1 ,\r8/t2/t0/s0/out_reg_n_2 ,\r8/t2/t0/s0/out_reg_n_3 ,\r8/t2/t0/s0/out_reg_n_4 ,\r8/t2/t0/s0/out_reg_n_5 ,\r8/t2/t0/s0/out_reg_n_6 ,\r8/t2/t0/s0/out_reg_n_7 ,\r8/t2/t0/p_0_in }),
        .DOBDO({\r8/t2/t0/s0/out_reg_n_16 ,\r8/t2/t0/s0/out_reg_n_17 ,\r8/t2/t0/s0/out_reg_n_18 ,\r8/t2/t0/s0/out_reg_n_19 ,\r8/t2/t0/s0/out_reg_n_20 ,\r8/t2/t0/s0/out_reg_n_21 ,\r8/t2/t0/s0/out_reg_n_22 ,\r8/t2/t0/s0/out_reg_n_23 ,\r8/t2/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r8/t2/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[63:56],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[55:48],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r8/t2/t0/s4/out_reg_n_0 ,\r8/t2/t0/s4/out_reg_n_1 ,\r8/t2/t0/s4/out_reg_n_2 ,\r8/t2/t0/s4/out_reg_n_3 ,\r8/t2/t0/s4/out_reg_n_4 ,\r8/t2/t0/s4/out_reg_n_5 ,\r8/t2/t0/s4/out_reg_n_6 ,\r8/t2/t0/s4/out_reg_n_7 ,\r8/t2/t0/p_1_in }),
        .DOBDO({\r8/t2/t0/s4/out_reg_n_16 ,\r8/t2/t0/s4/out_reg_n_17 ,\r8/t2/t0/s4/out_reg_n_18 ,\r8/t2/t0/s4/out_reg_n_19 ,\r8/t2/t0/s4/out_reg_n_20 ,\r8/t2/t0/s4/out_reg_n_21 ,\r8/t2/t0/s4/out_reg_n_22 ,\r8/t2/t0/s4/out_reg_n_23 ,\r8/t2/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r8/t2/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[47:40],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[39:32],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r8/t2/t2/s0/out_reg_n_0 ,\r8/t2/t2/s0/out_reg_n_1 ,\r8/t2/t2/s0/out_reg_n_2 ,\r8/t2/t2/s0/out_reg_n_3 ,\r8/t2/t2/s0/out_reg_n_4 ,\r8/t2/t2/s0/out_reg_n_5 ,\r8/t2/t2/s0/out_reg_n_6 ,\r8/t2/t2/s0/out_reg_n_7 ,\r8/t2/t2/p_0_in }),
        .DOBDO({\r8/t2/t2/s0/out_reg_n_16 ,\r8/t2/t2/s0/out_reg_n_17 ,\r8/t2/t2/s0/out_reg_n_18 ,\r8/t2/t2/s0/out_reg_n_19 ,\r8/t2/t2/s0/out_reg_n_20 ,\r8/t2/t2/s0/out_reg_n_21 ,\r8/t2/t2/s0/out_reg_n_22 ,\r8/t2/t2/s0/out_reg_n_23 ,\r8/t2/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r8/t2/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[47:40],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[39:32],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r8/t2/t2/s4/out_reg_n_0 ,\r8/t2/t2/s4/out_reg_n_1 ,\r8/t2/t2/s4/out_reg_n_2 ,\r8/t2/t2/s4/out_reg_n_3 ,\r8/t2/t2/s4/out_reg_n_4 ,\r8/t2/t2/s4/out_reg_n_5 ,\r8/t2/t2/s4/out_reg_n_6 ,\r8/t2/t2/s4/out_reg_n_7 ,\r8/t2/t2/p_1_in }),
        .DOBDO({\r8/t2/t2/s4/out_reg_n_16 ,\r8/t2/t2/s4/out_reg_n_17 ,\r8/t2/t2/s4/out_reg_n_18 ,\r8/t2/t2/s4/out_reg_n_19 ,\r8/t2/t2/s4/out_reg_n_20 ,\r8/t2/t2/s4/out_reg_n_21 ,\r8/t2/t2/s4/out_reg_n_22 ,\r8/t2/t2/s4/out_reg_n_23 ,\r8/t2/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r8/t3/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r8/t3/t0/s0/out_reg_n_0 ,\r8/t3/t0/s0/out_reg_n_1 ,\r8/t3/t0/s0/out_reg_n_2 ,\r8/t3/t0/s0/out_reg_n_3 ,\r8/t3/t0/s0/out_reg_n_4 ,\r8/t3/t0/s0/out_reg_n_5 ,\r8/t3/t0/s0/out_reg_n_6 ,\r8/t3/t0/s0/out_reg_n_7 ,\r8/t3/t0/p_0_in }),
        .DOBDO({\r8/t3/t0/s0/out_reg_n_16 ,\r8/t3/t0/s0/out_reg_n_17 ,\r8/t3/t0/s0/out_reg_n_18 ,\r8/t3/t0/s0/out_reg_n_19 ,\r8/t3/t0/s0/out_reg_n_20 ,\r8/t3/t0/s0/out_reg_n_21 ,\r8/t3/t0/s0/out_reg_n_22 ,\r8/t3/t0/s0/out_reg_n_23 ,\r8/t3/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r8/t3/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r8/t3/t0/s4/out_reg_n_0 ,\r8/t3/t0/s4/out_reg_n_1 ,\r8/t3/t0/s4/out_reg_n_2 ,\r8/t3/t0/s4/out_reg_n_3 ,\r8/t3/t0/s4/out_reg_n_4 ,\r8/t3/t0/s4/out_reg_n_5 ,\r8/t3/t0/s4/out_reg_n_6 ,\r8/t3/t0/s4/out_reg_n_7 ,\r8/t3/t0/p_1_in }),
        .DOBDO({\r8/t3/t0/s4/out_reg_n_16 ,\r8/t3/t0/s4/out_reg_n_17 ,\r8/t3/t0/s4/out_reg_n_18 ,\r8/t3/t0/s4/out_reg_n_19 ,\r8/t3/t0/s4/out_reg_n_20 ,\r8/t3/t0/s4/out_reg_n_21 ,\r8/t3/t0/s4/out_reg_n_22 ,\r8/t3/t0/s4/out_reg_n_23 ,\r8/t3/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r8/t3/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r8/t3/t2/s0/out_reg_n_0 ,\r8/t3/t2/s0/out_reg_n_1 ,\r8/t3/t2/s0/out_reg_n_2 ,\r8/t3/t2/s0/out_reg_n_3 ,\r8/t3/t2/s0/out_reg_n_4 ,\r8/t3/t2/s0/out_reg_n_5 ,\r8/t3/t2/s0/out_reg_n_6 ,\r8/t3/t2/s0/out_reg_n_7 ,\r8/t3/t2/p_0_in }),
        .DOBDO({\r8/t3/t2/s0/out_reg_n_16 ,\r8/t3/t2/s0/out_reg_n_17 ,\r8/t3/t2/s0/out_reg_n_18 ,\r8/t3/t2/s0/out_reg_n_19 ,\r8/t3/t2/s0/out_reg_n_20 ,\r8/t3/t2/s0/out_reg_n_21 ,\r8/t3/t2/s0/out_reg_n_22 ,\r8/t3/t2/s0/out_reg_n_23 ,\r8/t3/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r8/t3/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s7[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r8/t3/t2/s4/out_reg_n_0 ,\r8/t3/t2/s4/out_reg_n_1 ,\r8/t3/t2/s4/out_reg_n_2 ,\r8/t3/t2/s4/out_reg_n_3 ,\r8/t3/t2/s4/out_reg_n_4 ,\r8/t3/t2/s4/out_reg_n_5 ,\r8/t3/t2/s4/out_reg_n_6 ,\r8/t3/t2/s4/out_reg_n_7 ,\r8/t3/t2/p_1_in }),
        .DOBDO({\r8/t3/t2/s4/out_reg_n_16 ,\r8/t3/t2/s4/out_reg_n_17 ,\r8/t3/t2/s4/out_reg_n_18 ,\r8/t3/t2/s4/out_reg_n_19 ,\r8/t3/t2/s4/out_reg_n_20 ,\r8/t3/t2/s4/out_reg_n_21 ,\r8/t3/t2/s4/out_reg_n_22 ,\r8/t3/t2/s4/out_reg_n_23 ,\r8/t3/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [0]),
        .Q(s9[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[100] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [100]),
        .Q(s9[100]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[101] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [101]),
        .Q(s9[101]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[102] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [102]),
        .Q(s9[102]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[103] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [103]),
        .Q(s9[103]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[104] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [104]),
        .Q(s9[104]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[105] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [105]),
        .Q(s9[105]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[106] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [106]),
        .Q(s9[106]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[107] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [107]),
        .Q(s9[107]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[108] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [108]),
        .Q(s9[108]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[109] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [109]),
        .Q(s9[109]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [10]),
        .Q(s9[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[110] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [110]),
        .Q(s9[110]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[111] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [111]),
        .Q(s9[111]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[112] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [112]),
        .Q(s9[112]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[113] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [113]),
        .Q(s9[113]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[114] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [114]),
        .Q(s9[114]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[115] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [115]),
        .Q(s9[115]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[116] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [116]),
        .Q(s9[116]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[117] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [117]),
        .Q(s9[117]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[118] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [118]),
        .Q(s9[118]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[119] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [119]),
        .Q(s9[119]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [11]),
        .Q(s9[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[120] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [120]),
        .Q(s9[120]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[121] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [121]),
        .Q(s9[121]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[122] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [122]),
        .Q(s9[122]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[123] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [123]),
        .Q(s9[123]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[124] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [124]),
        .Q(s9[124]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[125] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [125]),
        .Q(s9[125]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[126] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [126]),
        .Q(s9[126]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[127] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [127]),
        .Q(s9[127]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [12]),
        .Q(s9[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [13]),
        .Q(s9[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [14]),
        .Q(s9[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [15]),
        .Q(s9[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [16]),
        .Q(s9[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [17]),
        .Q(s9[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [18]),
        .Q(s9[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [19]),
        .Q(s9[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [1]),
        .Q(s9[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [20]),
        .Q(s9[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [21]),
        .Q(s9[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [22]),
        .Q(s9[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [23]),
        .Q(s9[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [24]),
        .Q(s9[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [25]),
        .Q(s9[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [26]),
        .Q(s9[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [27]),
        .Q(s9[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [28]),
        .Q(s9[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [29]),
        .Q(s9[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [2]),
        .Q(s9[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [30]),
        .Q(s9[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [31]),
        .Q(s9[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [32]),
        .Q(s9[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [33]),
        .Q(s9[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [34]),
        .Q(s9[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [35]),
        .Q(s9[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [36]),
        .Q(s9[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [37]),
        .Q(s9[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [38]),
        .Q(s9[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [39]),
        .Q(s9[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [3]),
        .Q(s9[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [40]),
        .Q(s9[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [41]),
        .Q(s9[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [42]),
        .Q(s9[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [43]),
        .Q(s9[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [44]),
        .Q(s9[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [45]),
        .Q(s9[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [46]),
        .Q(s9[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [47]),
        .Q(s9[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [48]),
        .Q(s9[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [49]),
        .Q(s9[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [4]),
        .Q(s9[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [50]),
        .Q(s9[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [51]),
        .Q(s9[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [52]),
        .Q(s9[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [53]),
        .Q(s9[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [54]),
        .Q(s9[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [55]),
        .Q(s9[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [56]),
        .Q(s9[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [57]),
        .Q(s9[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [58]),
        .Q(s9[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [59]),
        .Q(s9[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [5]),
        .Q(s9[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [60]),
        .Q(s9[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [61]),
        .Q(s9[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [62]),
        .Q(s9[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [63]),
        .Q(s9[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[64] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [64]),
        .Q(s9[64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[65] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [65]),
        .Q(s9[65]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[66] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [66]),
        .Q(s9[66]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[67] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [67]),
        .Q(s9[67]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[68] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [68]),
        .Q(s9[68]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[69] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [69]),
        .Q(s9[69]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [6]),
        .Q(s9[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[70] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [70]),
        .Q(s9[70]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[71] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [71]),
        .Q(s9[71]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[72] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [72]),
        .Q(s9[72]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[73] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [73]),
        .Q(s9[73]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[74] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [74]),
        .Q(s9[74]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[75] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [75]),
        .Q(s9[75]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[76] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [76]),
        .Q(s9[76]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[77] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [77]),
        .Q(s9[77]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[78] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [78]),
        .Q(s9[78]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[79] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [79]),
        .Q(s9[79]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [7]),
        .Q(s9[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[80] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [80]),
        .Q(s9[80]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[81] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [81]),
        .Q(s9[81]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[82] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [82]),
        .Q(s9[82]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[83] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [83]),
        .Q(s9[83]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[84] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [84]),
        .Q(s9[84]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[85] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [85]),
        .Q(s9[85]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[86] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [86]),
        .Q(s9[86]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[87] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [87]),
        .Q(s9[87]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[88] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [88]),
        .Q(s9[88]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[89] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [89]),
        .Q(s9[89]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [8]),
        .Q(s9[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[90] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [90]),
        .Q(s9[90]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[91] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [91]),
        .Q(s9[91]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[92] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [92]),
        .Q(s9[92]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[93] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [93]),
        .Q(s9[93]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[94] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [94]),
        .Q(s9[94]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[95] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [95]),
        .Q(s9[95]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[96] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [96]),
        .Q(s9[96]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[97] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [97]),
        .Q(s9[97]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[98] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [98]),
        .Q(s9[98]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[99] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [99]),
        .Q(s9[99]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r9/state_out_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r9/p_0_out [9]),
        .Q(s9[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r9/t0/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[127:120],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[119:112],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r9/t0/t0/s0/out_reg_n_0 ,\r9/t0/t0/s0/out_reg_n_1 ,\r9/t0/t0/s0/out_reg_n_2 ,\r9/t0/t0/s0/out_reg_n_3 ,\r9/t0/t0/s0/out_reg_n_4 ,\r9/t0/t0/s0/out_reg_n_5 ,\r9/t0/t0/s0/out_reg_n_6 ,\r9/t0/t0/s0/out_reg_n_7 ,\r9/t0/t0/p_0_in }),
        .DOBDO({\r9/t0/t0/s0/out_reg_n_16 ,\r9/t0/t0/s0/out_reg_n_17 ,\r9/t0/t0/s0/out_reg_n_18 ,\r9/t0/t0/s0/out_reg_n_19 ,\r9/t0/t0/s0/out_reg_n_20 ,\r9/t0/t0/s0/out_reg_n_21 ,\r9/t0/t0/s0/out_reg_n_22 ,\r9/t0/t0/s0/out_reg_n_23 ,\r9/t0/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r9/t0/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[127:120],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[119:112],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r9/t0/t0/s4/out_reg_n_0 ,\r9/t0/t0/s4/out_reg_n_1 ,\r9/t0/t0/s4/out_reg_n_2 ,\r9/t0/t0/s4/out_reg_n_3 ,\r9/t0/t0/s4/out_reg_n_4 ,\r9/t0/t0/s4/out_reg_n_5 ,\r9/t0/t0/s4/out_reg_n_6 ,\r9/t0/t0/s4/out_reg_n_7 ,\r9/t0/t0/p_1_in }),
        .DOBDO({\r9/t0/t0/s4/out_reg_n_16 ,\r9/t0/t0/s4/out_reg_n_17 ,\r9/t0/t0/s4/out_reg_n_18 ,\r9/t0/t0/s4/out_reg_n_19 ,\r9/t0/t0/s4/out_reg_n_20 ,\r9/t0/t0/s4/out_reg_n_21 ,\r9/t0/t0/s4/out_reg_n_22 ,\r9/t0/t0/s4/out_reg_n_23 ,\r9/t0/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r9/t0/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[111:104],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[103:96],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r9/t0/t2/s0/out_reg_n_0 ,\r9/t0/t2/s0/out_reg_n_1 ,\r9/t0/t2/s0/out_reg_n_2 ,\r9/t0/t2/s0/out_reg_n_3 ,\r9/t0/t2/s0/out_reg_n_4 ,\r9/t0/t2/s0/out_reg_n_5 ,\r9/t0/t2/s0/out_reg_n_6 ,\r9/t0/t2/s0/out_reg_n_7 ,\r9/t0/t2/p_0_in }),
        .DOBDO({\r9/t0/t2/s0/out_reg_n_16 ,\r9/t0/t2/s0/out_reg_n_17 ,\r9/t0/t2/s0/out_reg_n_18 ,\r9/t0/t2/s0/out_reg_n_19 ,\r9/t0/t2/s0/out_reg_n_20 ,\r9/t0/t2/s0/out_reg_n_21 ,\r9/t0/t2/s0/out_reg_n_22 ,\r9/t0/t2/s0/out_reg_n_23 ,\r9/t0/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t0/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r9/t0/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[111:104],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[103:96],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r9/t0/t2/s4/out_reg_n_0 ,\r9/t0/t2/s4/out_reg_n_1 ,\r9/t0/t2/s4/out_reg_n_2 ,\r9/t0/t2/s4/out_reg_n_3 ,\r9/t0/t2/s4/out_reg_n_4 ,\r9/t0/t2/s4/out_reg_n_5 ,\r9/t0/t2/s4/out_reg_n_6 ,\r9/t0/t2/s4/out_reg_n_7 ,\r9/t0/t2/p_1_in }),
        .DOBDO({\r9/t0/t2/s4/out_reg_n_16 ,\r9/t0/t2/s4/out_reg_n_17 ,\r9/t0/t2/s4/out_reg_n_18 ,\r9/t0/t2/s4/out_reg_n_19 ,\r9/t0/t2/s4/out_reg_n_20 ,\r9/t0/t2/s4/out_reg_n_21 ,\r9/t0/t2/s4/out_reg_n_22 ,\r9/t0/t2/s4/out_reg_n_23 ,\r9/t0/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r9/t1/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[95:88],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[87:80],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r9/t1/t0/s0/out_reg_n_0 ,\r9/t1/t0/s0/out_reg_n_1 ,\r9/t1/t0/s0/out_reg_n_2 ,\r9/t1/t0/s0/out_reg_n_3 ,\r9/t1/t0/s0/out_reg_n_4 ,\r9/t1/t0/s0/out_reg_n_5 ,\r9/t1/t0/s0/out_reg_n_6 ,\r9/t1/t0/s0/out_reg_n_7 ,\r9/t1/t0/p_0_in }),
        .DOBDO({\r9/t1/t0/s0/out_reg_n_16 ,\r9/t1/t0/s0/out_reg_n_17 ,\r9/t1/t0/s0/out_reg_n_18 ,\r9/t1/t0/s0/out_reg_n_19 ,\r9/t1/t0/s0/out_reg_n_20 ,\r9/t1/t0/s0/out_reg_n_21 ,\r9/t1/t0/s0/out_reg_n_22 ,\r9/t1/t0/s0/out_reg_n_23 ,\r9/t1/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r9/t1/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[95:88],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[87:80],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r9/t1/t0/s4/out_reg_n_0 ,\r9/t1/t0/s4/out_reg_n_1 ,\r9/t1/t0/s4/out_reg_n_2 ,\r9/t1/t0/s4/out_reg_n_3 ,\r9/t1/t0/s4/out_reg_n_4 ,\r9/t1/t0/s4/out_reg_n_5 ,\r9/t1/t0/s4/out_reg_n_6 ,\r9/t1/t0/s4/out_reg_n_7 ,\r9/t1/t0/p_1_in }),
        .DOBDO({\r9/t1/t0/s4/out_reg_n_16 ,\r9/t1/t0/s4/out_reg_n_17 ,\r9/t1/t0/s4/out_reg_n_18 ,\r9/t1/t0/s4/out_reg_n_19 ,\r9/t1/t0/s4/out_reg_n_20 ,\r9/t1/t0/s4/out_reg_n_21 ,\r9/t1/t0/s4/out_reg_n_22 ,\r9/t1/t0/s4/out_reg_n_23 ,\r9/t1/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r9/t1/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[79:72],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[71:64],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r9/t1/t2/s0/out_reg_n_0 ,\r9/t1/t2/s0/out_reg_n_1 ,\r9/t1/t2/s0/out_reg_n_2 ,\r9/t1/t2/s0/out_reg_n_3 ,\r9/t1/t2/s0/out_reg_n_4 ,\r9/t1/t2/s0/out_reg_n_5 ,\r9/t1/t2/s0/out_reg_n_6 ,\r9/t1/t2/s0/out_reg_n_7 ,\r9/t1/t2/p_0_in }),
        .DOBDO({\r9/t1/t2/s0/out_reg_n_16 ,\r9/t1/t2/s0/out_reg_n_17 ,\r9/t1/t2/s0/out_reg_n_18 ,\r9/t1/t2/s0/out_reg_n_19 ,\r9/t1/t2/s0/out_reg_n_20 ,\r9/t1/t2/s0/out_reg_n_21 ,\r9/t1/t2/s0/out_reg_n_22 ,\r9/t1/t2/s0/out_reg_n_23 ,\r9/t1/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t1/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r9/t1/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[79:72],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[71:64],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r9/t1/t2/s4/out_reg_n_0 ,\r9/t1/t2/s4/out_reg_n_1 ,\r9/t1/t2/s4/out_reg_n_2 ,\r9/t1/t2/s4/out_reg_n_3 ,\r9/t1/t2/s4/out_reg_n_4 ,\r9/t1/t2/s4/out_reg_n_5 ,\r9/t1/t2/s4/out_reg_n_6 ,\r9/t1/t2/s4/out_reg_n_7 ,\r9/t1/t2/p_1_in }),
        .DOBDO({\r9/t1/t2/s4/out_reg_n_16 ,\r9/t1/t2/s4/out_reg_n_17 ,\r9/t1/t2/s4/out_reg_n_18 ,\r9/t1/t2/s4/out_reg_n_19 ,\r9/t1/t2/s4/out_reg_n_20 ,\r9/t1/t2/s4/out_reg_n_21 ,\r9/t1/t2/s4/out_reg_n_22 ,\r9/t1/t2/s4/out_reg_n_23 ,\r9/t1/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r9/t2/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[63:56],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[55:48],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r9/t2/t0/s0/out_reg_n_0 ,\r9/t2/t0/s0/out_reg_n_1 ,\r9/t2/t0/s0/out_reg_n_2 ,\r9/t2/t0/s0/out_reg_n_3 ,\r9/t2/t0/s0/out_reg_n_4 ,\r9/t2/t0/s0/out_reg_n_5 ,\r9/t2/t0/s0/out_reg_n_6 ,\r9/t2/t0/s0/out_reg_n_7 ,\r9/t2/t0/p_0_in }),
        .DOBDO({\r9/t2/t0/s0/out_reg_n_16 ,\r9/t2/t0/s0/out_reg_n_17 ,\r9/t2/t0/s0/out_reg_n_18 ,\r9/t2/t0/s0/out_reg_n_19 ,\r9/t2/t0/s0/out_reg_n_20 ,\r9/t2/t0/s0/out_reg_n_21 ,\r9/t2/t0/s0/out_reg_n_22 ,\r9/t2/t0/s0/out_reg_n_23 ,\r9/t2/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r9/t2/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[63:56],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[55:48],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r9/t2/t0/s4/out_reg_n_0 ,\r9/t2/t0/s4/out_reg_n_1 ,\r9/t2/t0/s4/out_reg_n_2 ,\r9/t2/t0/s4/out_reg_n_3 ,\r9/t2/t0/s4/out_reg_n_4 ,\r9/t2/t0/s4/out_reg_n_5 ,\r9/t2/t0/s4/out_reg_n_6 ,\r9/t2/t0/s4/out_reg_n_7 ,\r9/t2/t0/p_1_in }),
        .DOBDO({\r9/t2/t0/s4/out_reg_n_16 ,\r9/t2/t0/s4/out_reg_n_17 ,\r9/t2/t0/s4/out_reg_n_18 ,\r9/t2/t0/s4/out_reg_n_19 ,\r9/t2/t0/s4/out_reg_n_20 ,\r9/t2/t0/s4/out_reg_n_21 ,\r9/t2/t0/s4/out_reg_n_22 ,\r9/t2/t0/s4/out_reg_n_23 ,\r9/t2/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r9/t2/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[47:40],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[39:32],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r9/t2/t2/s0/out_reg_n_0 ,\r9/t2/t2/s0/out_reg_n_1 ,\r9/t2/t2/s0/out_reg_n_2 ,\r9/t2/t2/s0/out_reg_n_3 ,\r9/t2/t2/s0/out_reg_n_4 ,\r9/t2/t2/s0/out_reg_n_5 ,\r9/t2/t2/s0/out_reg_n_6 ,\r9/t2/t2/s0/out_reg_n_7 ,\r9/t2/t2/p_0_in }),
        .DOBDO({\r9/t2/t2/s0/out_reg_n_16 ,\r9/t2/t2/s0/out_reg_n_17 ,\r9/t2/t2/s0/out_reg_n_18 ,\r9/t2/t2/s0/out_reg_n_19 ,\r9/t2/t2/s0/out_reg_n_20 ,\r9/t2/t2/s0/out_reg_n_21 ,\r9/t2/t2/s0/out_reg_n_22 ,\r9/t2/t2/s0/out_reg_n_23 ,\r9/t2/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t2/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r9/t2/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[47:40],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[39:32],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r9/t2/t2/s4/out_reg_n_0 ,\r9/t2/t2/s4/out_reg_n_1 ,\r9/t2/t2/s4/out_reg_n_2 ,\r9/t2/t2/s4/out_reg_n_3 ,\r9/t2/t2/s4/out_reg_n_4 ,\r9/t2/t2/s4/out_reg_n_5 ,\r9/t2/t2/s4/out_reg_n_6 ,\r9/t2/t2/s4/out_reg_n_7 ,\r9/t2/t2/p_1_in }),
        .DOBDO({\r9/t2/t2/s4/out_reg_n_16 ,\r9/t2/t2/s4/out_reg_n_17 ,\r9/t2/t2/s4/out_reg_n_18 ,\r9/t2/t2/s4/out_reg_n_19 ,\r9/t2/t2/s4/out_reg_n_20 ,\r9/t2/t2/s4/out_reg_n_21 ,\r9/t2/t2/s4/out_reg_n_22 ,\r9/t2/t2/s4/out_reg_n_23 ,\r9/t2/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t0/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r9/t3/t0/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r9/t3/t0/s0/out_reg_n_0 ,\r9/t3/t0/s0/out_reg_n_1 ,\r9/t3/t0/s0/out_reg_n_2 ,\r9/t3/t0/s0/out_reg_n_3 ,\r9/t3/t0/s0/out_reg_n_4 ,\r9/t3/t0/s0/out_reg_n_5 ,\r9/t3/t0/s0/out_reg_n_6 ,\r9/t3/t0/s0/out_reg_n_7 ,\r9/t3/t0/p_0_in }),
        .DOBDO({\r9/t3/t0/s0/out_reg_n_16 ,\r9/t3/t0/s0/out_reg_n_17 ,\r9/t3/t0/s0/out_reg_n_18 ,\r9/t3/t0/s0/out_reg_n_19 ,\r9/t3/t0/s0/out_reg_n_20 ,\r9/t3/t0/s0/out_reg_n_21 ,\r9/t3/t0/s0/out_reg_n_22 ,\r9/t3/t0/s0/out_reg_n_23 ,\r9/t3/t1/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t0/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r9/t3/t0/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r9/t3/t0/s4/out_reg_n_0 ,\r9/t3/t0/s4/out_reg_n_1 ,\r9/t3/t0/s4/out_reg_n_2 ,\r9/t3/t0/s4/out_reg_n_3 ,\r9/t3/t0/s4/out_reg_n_4 ,\r9/t3/t0/s4/out_reg_n_5 ,\r9/t3/t0/s4/out_reg_n_6 ,\r9/t3/t0/s4/out_reg_n_7 ,\r9/t3/t0/p_1_in }),
        .DOBDO({\r9/t3/t0/s4/out_reg_n_16 ,\r9/t3/t0/s4/out_reg_n_17 ,\r9/t3/t0/s4/out_reg_n_18 ,\r9/t3/t0/s4/out_reg_n_19 ,\r9/t3/t0/s4/out_reg_n_20 ,\r9/t3/t0/s4/out_reg_n_21 ,\r9/t3/t0/s4/out_reg_n_22 ,\r9/t3/t0/s4/out_reg_n_23 ,\r9/t3/t1/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t2/s0/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r9/t3/t2/s0/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r9/t3/t2/s0/out_reg_n_0 ,\r9/t3/t2/s0/out_reg_n_1 ,\r9/t3/t2/s0/out_reg_n_2 ,\r9/t3/t2/s0/out_reg_n_3 ,\r9/t3/t2/s0/out_reg_n_4 ,\r9/t3/t2/s0/out_reg_n_5 ,\r9/t3/t2/s0/out_reg_n_6 ,\r9/t3/t2/s0/out_reg_n_7 ,\r9/t3/t2/p_0_in }),
        .DOBDO({\r9/t3/t2/s0/out_reg_n_16 ,\r9/t3/t2/s0/out_reg_n_17 ,\r9/t3/t2/s0/out_reg_n_18 ,\r9/t3/t2/s0/out_reg_n_19 ,\r9/t3/t2/s0/out_reg_n_20 ,\r9/t3/t2/s0/out_reg_n_21 ,\r9/t3/t2/s0/out_reg_n_22 ,\r9/t3/t2/s0/out_reg_n_23 ,\r9/t3/t3/p_0_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "t3/t2/s4/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00EC004D00B500E7005600CE00020060009100DE00D600FF00F600EE00F800C6),
    .INIT_01(256'h009B00E4005300230045005F00B3004100FB008E00B200EF00FA0089001F008F),
    .INIT_02(256'h002A006200AB00E200F900D100510068008300F5007E006C004C003D00E10075),
    .INIT_03(256'h00EA007F004E00CD00DF001B0024000E002F000A00370030009D004600950008),
    .INIT_04(256'h0013005E00DD0052007D00B7007600A4005B00B400DC003600340058001D0012),
    .INIT_05(256'h008500B00098009400720067008D00D400B6007900E3004000C1000000B900A6),
    .INIT_06(256'h004B0025007800A000FE000400E9008A00110066009A008600ED004F00C500BB),
    .INIT_07(256'h00BF00FD00E50020004200AF0077006300F100700021003F00050080005D00A2),
    .INIT_08(256'h00E6003200BA00C8007A00FC00550093002E0088003500BE00C3002600180081),
    .INIT_09(256'h00AD001600BC00A70028006B00C7008C000B003B0054004400A3009E001900C0),
    .INIT_0A(256'h00F200D30031003900C4004300BD009F00B80048000C009200140074006400DB),
    .INIT_0B(256'h0010004700F400CA00CF00F300AC00D80049009C00B1000100DA006E008B00D5),
    .INIT_0C(256'h000F000D00610096003E00E800A100CB0097007300570038005C004A00F0006F),
    .INIT_0D(256'h0027003A00990017006900AE006A00C2001C00F70006009000CC0071007C00E0),
    .INIT_0E(256'h00A5005000AA008700C90015003C002D0033000700A900D20022002B00EB00D9),
    .INIT_0F(256'h002C006D00A8007B001E005A0029008200D0008400D70065001A000900590003),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \r9/t3/t2/s4/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s8[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\r9/t3/t2/s4/out_reg_n_0 ,\r9/t3/t2/s4/out_reg_n_1 ,\r9/t3/t2/s4/out_reg_n_2 ,\r9/t3/t2/s4/out_reg_n_3 ,\r9/t3/t2/s4/out_reg_n_4 ,\r9/t3/t2/s4/out_reg_n_5 ,\r9/t3/t2/s4/out_reg_n_6 ,\r9/t3/t2/s4/out_reg_n_7 ,\r9/t3/t2/p_1_in }),
        .DOBDO({\r9/t3/t2/s4/out_reg_n_16 ,\r9/t3/t2/s4/out_reg_n_17 ,\r9/t3/t2/s4/out_reg_n_18 ,\r9/t3/t2/s4/out_reg_n_19 ,\r9/t3/t2/s4/out_reg_n_20 ,\r9/t3/t2/s4/out_reg_n_21 ,\r9/t3/t2/s4/out_reg_n_22 ,\r9/t3/t2/s4/out_reg_n_23 ,\r9/t3/t3/p_1_in }),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_1/S_1/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \rf/S4_1/S_1/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s9[119:112],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s9[127:120],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\rf/S4_1/S_1/out_reg_n_0 ,\rf/S4_1/S_1/out_reg_n_1 ,\rf/S4_1/S_1/out_reg_n_2 ,\rf/S4_1/S_1/out_reg_n_3 ,\rf/S4_1/S_1/out_reg_n_4 ,\rf/S4_1/S_1/out_reg_n_5 ,\rf/S4_1/S_1/out_reg_n_6 ,\rf/S4_1/S_1/out_reg_n_7 ,\rf/p_0_in [23:16]}),
        .DOBDO({\rf/S4_1/S_1/out_reg_n_16 ,\rf/S4_1/S_1/out_reg_n_17 ,\rf/S4_1/S_1/out_reg_n_18 ,\rf/S4_1/S_1/out_reg_n_19 ,\rf/S4_1/S_1/out_reg_n_20 ,\rf/S4_1/S_1/out_reg_n_21 ,\rf/S4_1/S_1/out_reg_n_22 ,\rf/S4_1/S_1/out_reg_n_23 ,\rf/p_3_in [31:24]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_1/S_3/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \rf/S4_1/S_3/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s9[103:96],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s9[111:104],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\rf/S4_1/S_3/out_reg_n_0 ,\rf/S4_1/S_3/out_reg_n_1 ,\rf/S4_1/S_3/out_reg_n_2 ,\rf/S4_1/S_3/out_reg_n_3 ,\rf/S4_1/S_3/out_reg_n_4 ,\rf/S4_1/S_3/out_reg_n_5 ,\rf/S4_1/S_3/out_reg_n_6 ,\rf/S4_1/S_3/out_reg_n_7 ,\rf/p_2_in [7:0]}),
        .DOBDO({\rf/S4_1/S_3/out_reg_n_16 ,\rf/S4_1/S_3/out_reg_n_17 ,\rf/S4_1/S_3/out_reg_n_18 ,\rf/S4_1/S_3/out_reg_n_19 ,\rf/S4_1/S_3/out_reg_n_20 ,\rf/S4_1/S_3/out_reg_n_21 ,\rf/S4_1/S_3/out_reg_n_22 ,\rf/S4_1/S_3/out_reg_n_23 ,\rf/p_1_in [15:8]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_2/S_1/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \rf/S4_2/S_1/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s9[87:80],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s9[95:88],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\rf/S4_2/S_1/out_reg_n_0 ,\rf/S4_2/S_1/out_reg_n_1 ,\rf/S4_2/S_1/out_reg_n_2 ,\rf/S4_2/S_1/out_reg_n_3 ,\rf/S4_2/S_1/out_reg_n_4 ,\rf/S4_2/S_1/out_reg_n_5 ,\rf/S4_2/S_1/out_reg_n_6 ,\rf/S4_2/S_1/out_reg_n_7 ,\rf/p_3_in [23:16]}),
        .DOBDO({\rf/S4_2/S_1/out_reg_n_16 ,\rf/S4_2/S_1/out_reg_n_17 ,\rf/S4_2/S_1/out_reg_n_18 ,\rf/S4_2/S_1/out_reg_n_19 ,\rf/S4_2/S_1/out_reg_n_20 ,\rf/S4_2/S_1/out_reg_n_21 ,\rf/S4_2/S_1/out_reg_n_22 ,\rf/S4_2/S_1/out_reg_n_23 ,\rf/p_2_in [31:24]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_2/S_3/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \rf/S4_2/S_3/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s9[71:64],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s9[79:72],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\rf/S4_2/S_3/out_reg_n_0 ,\rf/S4_2/S_3/out_reg_n_1 ,\rf/S4_2/S_3/out_reg_n_2 ,\rf/S4_2/S_3/out_reg_n_3 ,\rf/S4_2/S_3/out_reg_n_4 ,\rf/S4_2/S_3/out_reg_n_5 ,\rf/S4_2/S_3/out_reg_n_6 ,\rf/S4_2/S_3/out_reg_n_7 ,\rf/p_1_in [7:0]}),
        .DOBDO({\rf/S4_2/S_3/out_reg_n_16 ,\rf/S4_2/S_3/out_reg_n_17 ,\rf/S4_2/S_3/out_reg_n_18 ,\rf/S4_2/S_3/out_reg_n_19 ,\rf/S4_2/S_3/out_reg_n_20 ,\rf/S4_2/S_3/out_reg_n_21 ,\rf/S4_2/S_3/out_reg_n_22 ,\rf/S4_2/S_3/out_reg_n_23 ,\rf/p_0_in [15:8]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_3/S_1/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \rf/S4_3/S_1/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s9[55:48],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s9[63:56],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\rf/S4_3/S_1/out_reg_n_0 ,\rf/S4_3/S_1/out_reg_n_1 ,\rf/S4_3/S_1/out_reg_n_2 ,\rf/S4_3/S_1/out_reg_n_3 ,\rf/S4_3/S_1/out_reg_n_4 ,\rf/S4_3/S_1/out_reg_n_5 ,\rf/S4_3/S_1/out_reg_n_6 ,\rf/S4_3/S_1/out_reg_n_7 ,\rf/p_2_in [23:16]}),
        .DOBDO({\rf/S4_3/S_1/out_reg_n_16 ,\rf/S4_3/S_1/out_reg_n_17 ,\rf/S4_3/S_1/out_reg_n_18 ,\rf/S4_3/S_1/out_reg_n_19 ,\rf/S4_3/S_1/out_reg_n_20 ,\rf/S4_3/S_1/out_reg_n_21 ,\rf/S4_3/S_1/out_reg_n_22 ,\rf/S4_3/S_1/out_reg_n_23 ,\rf/p_1_in [31:24]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_3/S_3/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \rf/S4_3/S_3/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s9[39:32],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s9[47:40],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\rf/S4_3/S_3/out_reg_n_0 ,\rf/S4_3/S_3/out_reg_n_1 ,\rf/S4_3/S_3/out_reg_n_2 ,\rf/S4_3/S_3/out_reg_n_3 ,\rf/S4_3/S_3/out_reg_n_4 ,\rf/S4_3/S_3/out_reg_n_5 ,\rf/S4_3/S_3/out_reg_n_6 ,\rf/S4_3/S_3/out_reg_n_7 ,\rf/p_0_in [7:0]}),
        .DOBDO({\rf/S4_3/S_3/out_reg_n_16 ,\rf/S4_3/S_3/out_reg_n_17 ,\rf/S4_3/S_3/out_reg_n_18 ,\rf/S4_3/S_3/out_reg_n_19 ,\rf/S4_3/S_3/out_reg_n_20 ,\rf/S4_3/S_3/out_reg_n_21 ,\rf/S4_3/S_3/out_reg_n_22 ,\rf/S4_3/S_3/out_reg_n_23 ,\rf/p_3_in [15:8]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_4/S_1/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \rf/S4_4/S_1/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s9[23:16],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s9[31:24],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\rf/S4_4/S_1/out_reg_n_0 ,\rf/S4_4/S_1/out_reg_n_1 ,\rf/S4_4/S_1/out_reg_n_2 ,\rf/S4_4/S_1/out_reg_n_3 ,\rf/S4_4/S_1/out_reg_n_4 ,\rf/S4_4/S_1/out_reg_n_5 ,\rf/S4_4/S_1/out_reg_n_6 ,\rf/S4_4/S_1/out_reg_n_7 ,\rf/p_1_in [23:16]}),
        .DOBDO({\rf/S4_4/S_1/out_reg_n_16 ,\rf/S4_4/S_1/out_reg_n_17 ,\rf/S4_4/S_1/out_reg_n_18 ,\rf/S4_4/S_1/out_reg_n_19 ,\rf/S4_4/S_1/out_reg_n_20 ,\rf/S4_4/S_1/out_reg_n_21 ,\rf/S4_4/S_1/out_reg_n_22 ,\rf/S4_4/S_1/out_reg_n_23 ,\rf/p_0_in [31:24]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "2048" *) 
  (* RTL_RAM_NAME = "S4_4/S_3/out" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h007600AB00D700FE002B00670001003000C5006F006B00F2007B0077007C0063),
    .INIT_01(256'h00C0007200A4009C00AF00A200D400AD00F00047005900FA007D00C9008200CA),
    .INIT_02(256'h0015003100D8007100F100E500A5003400CC00F7003F00360026009300FD00B7),
    .INIT_03(256'h007500B2002700EB00E2008000120007009A00050096001800C3002300C70004),
    .INIT_04(256'h0084002F00E3002900B300D6003B005200A0005A006E001B001A002C00830009),
    .INIT_05(256'h00CF0058004C004A003900BE00CB006A005B00B100FC002000ED000000D10053),
    .INIT_06(256'h00A8009F003C0050007F000200F9004500850033004D004300FB00AA00EF00D0),
    .INIT_07(256'h00D200F300FF0010002100DA00B600BC00F50038009D0092008F004000A30051),
    .INIT_08(256'h00730019005D0064003D007E00A700C4001700440097005F00EC0013000C00CD),
    .INIT_09(256'h00DB000B005E00DE001400B800EE004600880090002A002200DC004F00810060),
    .INIT_0A(256'h007900E400950091006200AC00D300C2005C002400060049000A003A003200E0),
    .INIT_0B(256'h000800AE007A006500EA00F40056006C00A9004E00D5008D006D003700C800E7),
    .INIT_0C(256'h008A008B00BD004B001F007400DD00E800C600B400A6001C002E0025007800BA),
    .INIT_0D(256'h009E001D00C1008600B9005700350061000E00F600030048006600B5003E0070),
    .INIT_0E(256'h00DF0028005500CE00E90087001E009B0094008E00D900690011009800F800E1),
    .INIT_0F(256'h001600BB005400B0000F002D009900410068004200E600BF000D008900A1008C),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \rf/S4_4/S_3/out_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,s9[7:0],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,s9[15:8],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\rf/S4_4/S_3/out_reg_n_0 ,\rf/S4_4/S_3/out_reg_n_1 ,\rf/S4_4/S_3/out_reg_n_2 ,\rf/S4_4/S_3/out_reg_n_3 ,\rf/S4_4/S_3/out_reg_n_4 ,\rf/S4_4/S_3/out_reg_n_5 ,\rf/S4_4/S_3/out_reg_n_6 ,\rf/S4_4/S_3/out_reg_n_7 ,\rf/p_3_in [7:0]}),
        .DOBDO({\rf/S4_4/S_3/out_reg_n_16 ,\rf/S4_4/S_3/out_reg_n_17 ,\rf/S4_4/S_3/out_reg_n_18 ,\rf/S4_4/S_3/out_reg_n_19 ,\rf/S4_4/S_3/out_reg_n_20 ,\rf/S4_4/S_3/out_reg_n_21 ,\rf/S4_4/S_3/out_reg_n_22 ,\rf/S4_4/S_3/out_reg_n_23 ,\rf/p_2_in [15:8]}),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\<const1>__0__0 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [0]),
        .Q(out[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[100] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [100]),
        .Q(out[100]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[101] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [101]),
        .Q(out[101]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[102] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [102]),
        .Q(out[102]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[103] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [103]),
        .Q(out[103]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[104] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [104]),
        .Q(out[104]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[105] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [105]),
        .Q(out[105]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[106] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [106]),
        .Q(out[106]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[107] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [107]),
        .Q(out[107]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[108] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [108]),
        .Q(out[108]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[109] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [109]),
        .Q(out[109]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [10]),
        .Q(out[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[110] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [110]),
        .Q(out[110]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[111] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [111]),
        .Q(out[111]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[112] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [112]),
        .Q(out[112]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[113] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [113]),
        .Q(out[113]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[114] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [114]),
        .Q(out[114]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[115] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [115]),
        .Q(out[115]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[116] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [116]),
        .Q(out[116]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[117] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [117]),
        .Q(out[117]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[118] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [118]),
        .Q(out[118]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[119] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [119]),
        .Q(out[119]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [11]),
        .Q(out[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[120] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [120]),
        .Q(out[120]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[121] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [121]),
        .Q(out[121]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[122] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [122]),
        .Q(out[122]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[123] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [123]),
        .Q(out[123]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[124] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [124]),
        .Q(out[124]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[125] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [125]),
        .Q(out[125]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[126] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [126]),
        .Q(out[126]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[127] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [127]),
        .Q(out[127]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [12]),
        .Q(out[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [13]),
        .Q(out[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [14]),
        .Q(out[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [15]),
        .Q(out[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [16]),
        .Q(out[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [17]),
        .Q(out[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [18]),
        .Q(out[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [19]),
        .Q(out[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [1]),
        .Q(out[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [20]),
        .Q(out[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [21]),
        .Q(out[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [22]),
        .Q(out[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [23]),
        .Q(out[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [24]),
        .Q(out[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [25]),
        .Q(out[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [26]),
        .Q(out[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [27]),
        .Q(out[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [28]),
        .Q(out[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [29]),
        .Q(out[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [2]),
        .Q(out[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [30]),
        .Q(out[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [31]),
        .Q(out[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [32]),
        .Q(out[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [33]),
        .Q(out[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [34]),
        .Q(out[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [35]),
        .Q(out[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [36]),
        .Q(out[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [37]),
        .Q(out[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [38]),
        .Q(out[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [39]),
        .Q(out[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [3]),
        .Q(out[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [40]),
        .Q(out[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [41]),
        .Q(out[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [42]),
        .Q(out[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [43]),
        .Q(out[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [44]),
        .Q(out[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [45]),
        .Q(out[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [46]),
        .Q(out[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [47]),
        .Q(out[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [48]),
        .Q(out[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [49]),
        .Q(out[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [4]),
        .Q(out[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [50]),
        .Q(out[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [51]),
        .Q(out[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [52]),
        .Q(out[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [53]),
        .Q(out[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [54]),
        .Q(out[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [55]),
        .Q(out[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [56]),
        .Q(out[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [57]),
        .Q(out[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [58]),
        .Q(out[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [59]),
        .Q(out[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [5]),
        .Q(out[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [60]),
        .Q(out[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [61]),
        .Q(out[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [62]),
        .Q(out[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [63]),
        .Q(out[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[64] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [64]),
        .Q(out[64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[65] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [65]),
        .Q(out[65]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[66] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [66]),
        .Q(out[66]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[67] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [67]),
        .Q(out[67]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[68] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [68]),
        .Q(out[68]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[69] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [69]),
        .Q(out[69]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [6]),
        .Q(out[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[70] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [70]),
        .Q(out[70]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[71] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [71]),
        .Q(out[71]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[72] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [72]),
        .Q(out[72]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[73] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [73]),
        .Q(out[73]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[74] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [74]),
        .Q(out[74]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[75] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [75]),
        .Q(out[75]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[76] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [76]),
        .Q(out[76]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[77] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [77]),
        .Q(out[77]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[78] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [78]),
        .Q(out[78]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[79] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [79]),
        .Q(out[79]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [7]),
        .Q(out[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[80] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [80]),
        .Q(out[80]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[81] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [81]),
        .Q(out[81]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[82] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [82]),
        .Q(out[82]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[83] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [83]),
        .Q(out[83]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[84] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [84]),
        .Q(out[84]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[85] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [85]),
        .Q(out[85]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[86] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [86]),
        .Q(out[86]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[87] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [87]),
        .Q(out[87]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[88] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [88]),
        .Q(out[88]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[89] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [89]),
        .Q(out[89]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [8]),
        .Q(out[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[90] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [90]),
        .Q(out[90]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[91] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [91]),
        .Q(out[91]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[92] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [92]),
        .Q(out[92]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[93] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [93]),
        .Q(out[93]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[94] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [94]),
        .Q(out[94]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[95] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [95]),
        .Q(out[95]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[96] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [96]),
        .Q(out[96]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[97] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [97]),
        .Q(out[97]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[98] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [98]),
        .Q(out[98]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[99] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [99]),
        .Q(out[99]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \rf/state_out_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rf/p_4_out [9]),
        .Q(out[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[0]_i_1 
       (.I0(state[0]),
        .I1(key[0]),
        .O(\s0[0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[100]_i_1 
       (.I0(state[100]),
        .I1(key[100]),
        .O(\s0[100]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[101]_i_1 
       (.I0(state[101]),
        .I1(key[101]),
        .O(\s0[101]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[102]_i_1 
       (.I0(state[102]),
        .I1(key[102]),
        .O(\s0[102]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[103]_i_1 
       (.I0(state[103]),
        .I1(key[103]),
        .O(\s0[103]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[104]_i_1 
       (.I0(state[104]),
        .I1(key[104]),
        .O(\s0[104]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[105]_i_1 
       (.I0(state[105]),
        .I1(key[105]),
        .O(\s0[105]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[106]_i_1 
       (.I0(state[106]),
        .I1(key[106]),
        .O(\s0[106]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[107]_i_1 
       (.I0(state[107]),
        .I1(key[107]),
        .O(\s0[107]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[108]_i_1 
       (.I0(state[108]),
        .I1(key[108]),
        .O(\s0[108]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[109]_i_1 
       (.I0(state[109]),
        .I1(key[109]),
        .O(\s0[109]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[10]_i_1 
       (.I0(state[10]),
        .I1(key[10]),
        .O(\s0[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[110]_i_1 
       (.I0(state[110]),
        .I1(key[110]),
        .O(\s0[110]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[111]_i_1 
       (.I0(state[111]),
        .I1(key[111]),
        .O(\s0[111]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[112]_i_1 
       (.I0(state[112]),
        .I1(key[112]),
        .O(\s0[112]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[113]_i_1 
       (.I0(state[113]),
        .I1(key[113]),
        .O(\s0[113]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[114]_i_1 
       (.I0(state[114]),
        .I1(key[114]),
        .O(\s0[114]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[115]_i_1 
       (.I0(state[115]),
        .I1(key[115]),
        .O(\s0[115]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[116]_i_1 
       (.I0(state[116]),
        .I1(key[116]),
        .O(\s0[116]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[117]_i_1 
       (.I0(state[117]),
        .I1(key[117]),
        .O(\s0[117]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[118]_i_1 
       (.I0(state[118]),
        .I1(key[118]),
        .O(\s0[118]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[119]_i_1 
       (.I0(state[119]),
        .I1(key[119]),
        .O(\s0[119]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[11]_i_1 
       (.I0(state[11]),
        .I1(key[11]),
        .O(\s0[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[120]_i_1 
       (.I0(state[120]),
        .I1(key[120]),
        .O(\s0[120]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[121]_i_1 
       (.I0(state[121]),
        .I1(key[121]),
        .O(\s0[121]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[122]_i_1 
       (.I0(state[122]),
        .I1(key[122]),
        .O(\s0[122]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[123]_i_1 
       (.I0(state[123]),
        .I1(key[123]),
        .O(\s0[123]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[124]_i_1 
       (.I0(state[124]),
        .I1(key[124]),
        .O(\s0[124]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[125]_i_1 
       (.I0(state[125]),
        .I1(key[125]),
        .O(\s0[125]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[126]_i_1 
       (.I0(state[126]),
        .I1(key[126]),
        .O(\s0[126]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[127]_i_1 
       (.I0(state[127]),
        .I1(key[127]),
        .O(\s0[127]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[12]_i_1 
       (.I0(state[12]),
        .I1(key[12]),
        .O(\s0[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[13]_i_1 
       (.I0(state[13]),
        .I1(key[13]),
        .O(\s0[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[14]_i_1 
       (.I0(state[14]),
        .I1(key[14]),
        .O(\s0[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[15]_i_1 
       (.I0(state[15]),
        .I1(key[15]),
        .O(\s0[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[16]_i_1 
       (.I0(state[16]),
        .I1(key[16]),
        .O(\s0[16]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[17]_i_1 
       (.I0(state[17]),
        .I1(key[17]),
        .O(\s0[17]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[18]_i_1 
       (.I0(state[18]),
        .I1(key[18]),
        .O(\s0[18]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[19]_i_1 
       (.I0(state[19]),
        .I1(key[19]),
        .O(\s0[19]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[1]_i_1 
       (.I0(state[1]),
        .I1(key[1]),
        .O(\s0[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[20]_i_1 
       (.I0(state[20]),
        .I1(key[20]),
        .O(\s0[20]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[21]_i_1 
       (.I0(state[21]),
        .I1(key[21]),
        .O(\s0[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[22]_i_1 
       (.I0(state[22]),
        .I1(key[22]),
        .O(\s0[22]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[23]_i_1 
       (.I0(state[23]),
        .I1(key[23]),
        .O(\s0[23]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[24]_i_1 
       (.I0(state[24]),
        .I1(key[24]),
        .O(\s0[24]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[25]_i_1 
       (.I0(state[25]),
        .I1(key[25]),
        .O(\s0[25]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[26]_i_1 
       (.I0(state[26]),
        .I1(key[26]),
        .O(\s0[26]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[27]_i_1 
       (.I0(state[27]),
        .I1(key[27]),
        .O(\s0[27]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[28]_i_1 
       (.I0(state[28]),
        .I1(key[28]),
        .O(\s0[28]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[29]_i_1 
       (.I0(state[29]),
        .I1(key[29]),
        .O(\s0[29]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[2]_i_1 
       (.I0(state[2]),
        .I1(key[2]),
        .O(\s0[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[30]_i_1 
       (.I0(state[30]),
        .I1(key[30]),
        .O(\s0[30]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[31]_i_1 
       (.I0(state[31]),
        .I1(key[31]),
        .O(\s0[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[32]_i_1 
       (.I0(state[32]),
        .I1(key[32]),
        .O(\s0[32]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[33]_i_1 
       (.I0(state[33]),
        .I1(key[33]),
        .O(\s0[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[34]_i_1 
       (.I0(state[34]),
        .I1(key[34]),
        .O(\s0[34]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[35]_i_1 
       (.I0(state[35]),
        .I1(key[35]),
        .O(\s0[35]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[36]_i_1 
       (.I0(state[36]),
        .I1(key[36]),
        .O(\s0[36]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[37]_i_1 
       (.I0(state[37]),
        .I1(key[37]),
        .O(\s0[37]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[38]_i_1 
       (.I0(state[38]),
        .I1(key[38]),
        .O(\s0[38]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[39]_i_1 
       (.I0(state[39]),
        .I1(key[39]),
        .O(\s0[39]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[3]_i_1 
       (.I0(state[3]),
        .I1(key[3]),
        .O(\s0[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[40]_i_1 
       (.I0(state[40]),
        .I1(key[40]),
        .O(\s0[40]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[41]_i_1 
       (.I0(state[41]),
        .I1(key[41]),
        .O(\s0[41]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[42]_i_1 
       (.I0(state[42]),
        .I1(key[42]),
        .O(\s0[42]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[43]_i_1 
       (.I0(state[43]),
        .I1(key[43]),
        .O(\s0[43]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[44]_i_1 
       (.I0(state[44]),
        .I1(key[44]),
        .O(\s0[44]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[45]_i_1 
       (.I0(state[45]),
        .I1(key[45]),
        .O(\s0[45]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[46]_i_1 
       (.I0(state[46]),
        .I1(key[46]),
        .O(\s0[46]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[47]_i_1 
       (.I0(state[47]),
        .I1(key[47]),
        .O(\s0[47]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[48]_i_1 
       (.I0(state[48]),
        .I1(key[48]),
        .O(\s0[48]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[49]_i_1 
       (.I0(state[49]),
        .I1(key[49]),
        .O(\s0[49]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[4]_i_1 
       (.I0(state[4]),
        .I1(key[4]),
        .O(\s0[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[50]_i_1 
       (.I0(state[50]),
        .I1(key[50]),
        .O(\s0[50]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[51]_i_1 
       (.I0(state[51]),
        .I1(key[51]),
        .O(\s0[51]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[52]_i_1 
       (.I0(state[52]),
        .I1(key[52]),
        .O(\s0[52]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[53]_i_1 
       (.I0(state[53]),
        .I1(key[53]),
        .O(\s0[53]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[54]_i_1 
       (.I0(state[54]),
        .I1(key[54]),
        .O(\s0[54]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[55]_i_1 
       (.I0(state[55]),
        .I1(key[55]),
        .O(\s0[55]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[56]_i_1 
       (.I0(state[56]),
        .I1(key[56]),
        .O(\s0[56]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[57]_i_1 
       (.I0(state[57]),
        .I1(key[57]),
        .O(\s0[57]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[58]_i_1 
       (.I0(state[58]),
        .I1(key[58]),
        .O(\s0[58]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[59]_i_1 
       (.I0(state[59]),
        .I1(key[59]),
        .O(\s0[59]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[5]_i_1 
       (.I0(state[5]),
        .I1(key[5]),
        .O(\s0[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[60]_i_1 
       (.I0(state[60]),
        .I1(key[60]),
        .O(\s0[60]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[61]_i_1 
       (.I0(state[61]),
        .I1(key[61]),
        .O(\s0[61]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[62]_i_1 
       (.I0(state[62]),
        .I1(key[62]),
        .O(\s0[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[63]_i_1 
       (.I0(state[63]),
        .I1(key[63]),
        .O(\s0[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[64]_i_1 
       (.I0(state[64]),
        .I1(key[64]),
        .O(\s0[64]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[65]_i_1 
       (.I0(state[65]),
        .I1(key[65]),
        .O(\s0[65]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[66]_i_1 
       (.I0(state[66]),
        .I1(key[66]),
        .O(\s0[66]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[67]_i_1 
       (.I0(state[67]),
        .I1(key[67]),
        .O(\s0[67]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[68]_i_1 
       (.I0(state[68]),
        .I1(key[68]),
        .O(\s0[68]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[69]_i_1 
       (.I0(state[69]),
        .I1(key[69]),
        .O(\s0[69]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[6]_i_1 
       (.I0(state[6]),
        .I1(key[6]),
        .O(\s0[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[70]_i_1 
       (.I0(state[70]),
        .I1(key[70]),
        .O(\s0[70]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[71]_i_1 
       (.I0(state[71]),
        .I1(key[71]),
        .O(\s0[71]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[72]_i_1 
       (.I0(state[72]),
        .I1(key[72]),
        .O(\s0[72]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[73]_i_1 
       (.I0(state[73]),
        .I1(key[73]),
        .O(\s0[73]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[74]_i_1 
       (.I0(state[74]),
        .I1(key[74]),
        .O(\s0[74]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[75]_i_1 
       (.I0(state[75]),
        .I1(key[75]),
        .O(\s0[75]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[76]_i_1 
       (.I0(state[76]),
        .I1(key[76]),
        .O(\s0[76]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[77]_i_1 
       (.I0(state[77]),
        .I1(key[77]),
        .O(\s0[77]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[78]_i_1 
       (.I0(state[78]),
        .I1(key[78]),
        .O(\s0[78]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[79]_i_1 
       (.I0(state[79]),
        .I1(key[79]),
        .O(\s0[79]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[7]_i_1 
       (.I0(state[7]),
        .I1(key[7]),
        .O(\s0[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[80]_i_1 
       (.I0(state[80]),
        .I1(key[80]),
        .O(\s0[80]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[81]_i_1 
       (.I0(state[81]),
        .I1(key[81]),
        .O(\s0[81]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[82]_i_1 
       (.I0(state[82]),
        .I1(key[82]),
        .O(\s0[82]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[83]_i_1 
       (.I0(state[83]),
        .I1(key[83]),
        .O(\s0[83]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[84]_i_1 
       (.I0(state[84]),
        .I1(key[84]),
        .O(\s0[84]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[85]_i_1 
       (.I0(state[85]),
        .I1(key[85]),
        .O(\s0[85]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[86]_i_1 
       (.I0(state[86]),
        .I1(key[86]),
        .O(\s0[86]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[87]_i_1 
       (.I0(state[87]),
        .I1(key[87]),
        .O(\s0[87]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[88]_i_1 
       (.I0(state[88]),
        .I1(key[88]),
        .O(\s0[88]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[89]_i_1 
       (.I0(state[89]),
        .I1(key[89]),
        .O(\s0[89]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[8]_i_1 
       (.I0(state[8]),
        .I1(key[8]),
        .O(\s0[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[90]_i_1 
       (.I0(state[90]),
        .I1(key[90]),
        .O(\s0[90]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[91]_i_1 
       (.I0(state[91]),
        .I1(key[91]),
        .O(\s0[91]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[92]_i_1 
       (.I0(state[92]),
        .I1(key[92]),
        .O(\s0[92]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[93]_i_1 
       (.I0(state[93]),
        .I1(key[93]),
        .O(\s0[93]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[94]_i_1 
       (.I0(state[94]),
        .I1(key[94]),
        .O(\s0[94]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[95]_i_1 
       (.I0(state[95]),
        .I1(key[95]),
        .O(\s0[95]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[96]_i_1 
       (.I0(state[96]),
        .I1(key[96]),
        .O(\s0[96]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[97]_i_1 
       (.I0(state[97]),
        .I1(key[97]),
        .O(\s0[97]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[98]_i_1 
       (.I0(state[98]),
        .I1(key[98]),
        .O(\s0[98]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[99]_i_1 
       (.I0(state[99]),
        .I1(key[99]),
        .O(\s0[99]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \s0[9]_i_1 
       (.I0(state[9]),
        .I1(key[9]),
        .O(\s0[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[0]_i_1_n_0 ),
        .Q(s0[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[100] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[100]_i_1_n_0 ),
        .Q(s0[100]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[101] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[101]_i_1_n_0 ),
        .Q(s0[101]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[102] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[102]_i_1_n_0 ),
        .Q(s0[102]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[103] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[103]_i_1_n_0 ),
        .Q(s0[103]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[104] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[104]_i_1_n_0 ),
        .Q(s0[104]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[105] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[105]_i_1_n_0 ),
        .Q(s0[105]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[106] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[106]_i_1_n_0 ),
        .Q(s0[106]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[107] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[107]_i_1_n_0 ),
        .Q(s0[107]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[108] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[108]_i_1_n_0 ),
        .Q(s0[108]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[109] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[109]_i_1_n_0 ),
        .Q(s0[109]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[10]_i_1_n_0 ),
        .Q(s0[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[110] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[110]_i_1_n_0 ),
        .Q(s0[110]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[111] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[111]_i_1_n_0 ),
        .Q(s0[111]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[112] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[112]_i_1_n_0 ),
        .Q(s0[112]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[113] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[113]_i_1_n_0 ),
        .Q(s0[113]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[114] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[114]_i_1_n_0 ),
        .Q(s0[114]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[115] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[115]_i_1_n_0 ),
        .Q(s0[115]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[116] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[116]_i_1_n_0 ),
        .Q(s0[116]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[117] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[117]_i_1_n_0 ),
        .Q(s0[117]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[118] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[118]_i_1_n_0 ),
        .Q(s0[118]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[119] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[119]_i_1_n_0 ),
        .Q(s0[119]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[11]_i_1_n_0 ),
        .Q(s0[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[120] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[120]_i_1_n_0 ),
        .Q(s0[120]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[121] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[121]_i_1_n_0 ),
        .Q(s0[121]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[122] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[122]_i_1_n_0 ),
        .Q(s0[122]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[123] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[123]_i_1_n_0 ),
        .Q(s0[123]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[124] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[124]_i_1_n_0 ),
        .Q(s0[124]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[125] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[125]_i_1_n_0 ),
        .Q(s0[125]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[126] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[126]_i_1_n_0 ),
        .Q(s0[126]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[127] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[127]_i_1_n_0 ),
        .Q(s0[127]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[12]_i_1_n_0 ),
        .Q(s0[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[13]_i_1_n_0 ),
        .Q(s0[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[14]_i_1_n_0 ),
        .Q(s0[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[15]_i_1_n_0 ),
        .Q(s0[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[16]_i_1_n_0 ),
        .Q(s0[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[17]_i_1_n_0 ),
        .Q(s0[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[18]_i_1_n_0 ),
        .Q(s0[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[19]_i_1_n_0 ),
        .Q(s0[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[1]_i_1_n_0 ),
        .Q(s0[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[20]_i_1_n_0 ),
        .Q(s0[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[21]_i_1_n_0 ),
        .Q(s0[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[22]_i_1_n_0 ),
        .Q(s0[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[23]_i_1_n_0 ),
        .Q(s0[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[24]_i_1_n_0 ),
        .Q(s0[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[25]_i_1_n_0 ),
        .Q(s0[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[26]_i_1_n_0 ),
        .Q(s0[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[27]_i_1_n_0 ),
        .Q(s0[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[28]_i_1_n_0 ),
        .Q(s0[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[29]_i_1_n_0 ),
        .Q(s0[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[2]_i_1_n_0 ),
        .Q(s0[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[30]_i_1_n_0 ),
        .Q(s0[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[31]_i_1_n_0 ),
        .Q(s0[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[32]_i_1_n_0 ),
        .Q(s0[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[33]_i_1_n_0 ),
        .Q(s0[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[34]_i_1_n_0 ),
        .Q(s0[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[35]_i_1_n_0 ),
        .Q(s0[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[36]_i_1_n_0 ),
        .Q(s0[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[37]_i_1_n_0 ),
        .Q(s0[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[38]_i_1_n_0 ),
        .Q(s0[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[39]_i_1_n_0 ),
        .Q(s0[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[3]_i_1_n_0 ),
        .Q(s0[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[40]_i_1_n_0 ),
        .Q(s0[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[41]_i_1_n_0 ),
        .Q(s0[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[42]_i_1_n_0 ),
        .Q(s0[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[43]_i_1_n_0 ),
        .Q(s0[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[44]_i_1_n_0 ),
        .Q(s0[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[45]_i_1_n_0 ),
        .Q(s0[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[46]_i_1_n_0 ),
        .Q(s0[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[47]_i_1_n_0 ),
        .Q(s0[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[48]_i_1_n_0 ),
        .Q(s0[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[49]_i_1_n_0 ),
        .Q(s0[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[4]_i_1_n_0 ),
        .Q(s0[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[50]_i_1_n_0 ),
        .Q(s0[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[51]_i_1_n_0 ),
        .Q(s0[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[52]_i_1_n_0 ),
        .Q(s0[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[53]_i_1_n_0 ),
        .Q(s0[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[54]_i_1_n_0 ),
        .Q(s0[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[55]_i_1_n_0 ),
        .Q(s0[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[56]_i_1_n_0 ),
        .Q(s0[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[57]_i_1_n_0 ),
        .Q(s0[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[58]_i_1_n_0 ),
        .Q(s0[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[59]_i_1_n_0 ),
        .Q(s0[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[5]_i_1_n_0 ),
        .Q(s0[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[60]_i_1_n_0 ),
        .Q(s0[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[61]_i_1_n_0 ),
        .Q(s0[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[62]_i_1_n_0 ),
        .Q(s0[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[63]_i_1_n_0 ),
        .Q(s0[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[64] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[64]_i_1_n_0 ),
        .Q(s0[64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[65] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[65]_i_1_n_0 ),
        .Q(s0[65]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[66] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[66]_i_1_n_0 ),
        .Q(s0[66]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[67] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[67]_i_1_n_0 ),
        .Q(s0[67]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[68] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[68]_i_1_n_0 ),
        .Q(s0[68]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[69] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[69]_i_1_n_0 ),
        .Q(s0[69]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[6]_i_1_n_0 ),
        .Q(s0[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[70] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[70]_i_1_n_0 ),
        .Q(s0[70]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[71] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[71]_i_1_n_0 ),
        .Q(s0[71]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[72] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[72]_i_1_n_0 ),
        .Q(s0[72]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[73] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[73]_i_1_n_0 ),
        .Q(s0[73]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[74] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[74]_i_1_n_0 ),
        .Q(s0[74]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[75] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[75]_i_1_n_0 ),
        .Q(s0[75]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[76] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[76]_i_1_n_0 ),
        .Q(s0[76]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[77] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[77]_i_1_n_0 ),
        .Q(s0[77]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[78] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[78]_i_1_n_0 ),
        .Q(s0[78]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[79] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[79]_i_1_n_0 ),
        .Q(s0[79]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[7]_i_1_n_0 ),
        .Q(s0[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[80] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[80]_i_1_n_0 ),
        .Q(s0[80]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[81] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[81]_i_1_n_0 ),
        .Q(s0[81]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[82] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[82]_i_1_n_0 ),
        .Q(s0[82]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[83] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[83]_i_1_n_0 ),
        .Q(s0[83]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[84] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[84]_i_1_n_0 ),
        .Q(s0[84]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[85] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[85]_i_1_n_0 ),
        .Q(s0[85]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[86] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[86]_i_1_n_0 ),
        .Q(s0[86]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[87] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[87]_i_1_n_0 ),
        .Q(s0[87]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[88] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[88]_i_1_n_0 ),
        .Q(s0[88]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[89] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[89]_i_1_n_0 ),
        .Q(s0[89]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[8]_i_1_n_0 ),
        .Q(s0[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[90] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[90]_i_1_n_0 ),
        .Q(s0[90]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[91] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[91]_i_1_n_0 ),
        .Q(s0[91]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[92] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[92]_i_1_n_0 ),
        .Q(s0[92]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[93] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[93]_i_1_n_0 ),
        .Q(s0[93]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[94] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[94]_i_1_n_0 ),
        .Q(s0[94]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[95] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[95]_i_1_n_0 ),
        .Q(s0[95]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[96] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[96]_i_1_n_0 ),
        .Q(s0[96]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[97] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[97]_i_1_n_0 ),
        .Q(s0[97]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[98] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[98]_i_1_n_0 ),
        .Q(s0[98]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[99] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[99]_i_1_n_0 ),
        .Q(s0[99]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \s0_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\s0[9]_i_1_n_0 ),
        .Q(s0[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[0]_i_1 
       (.I0(\r1/t0/t1/p_0_in [0]),
        .I1(\r1/t2/t3/p_1_in [0]),
        .I2(\r1/t1/t2/p_0_in [0]),
        .I3(k0b[0]),
        .I4(\r1/t3/t0/p_1_in [0]),
        .I5(\r1/t3/t0/p_0_in [0]),
        .O(\r1/p_0_out [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[0]_i_1__0 
       (.I0(\r2/t0/t1/p_0_in [0]),
        .I1(\r2/t2/t3/p_1_in [0]),
        .I2(\r2/t1/t2/p_0_in [0]),
        .I3(k1b[0]),
        .I4(\r2/t3/t0/p_1_in [0]),
        .I5(\r2/t3/t0/p_0_in [0]),
        .O(\r2/p_0_out [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[0]_i_1__1 
       (.I0(\r3/t0/t1/p_0_in [0]),
        .I1(\r3/t2/t3/p_1_in [0]),
        .I2(\r3/t1/t2/p_0_in [0]),
        .I3(k2b[0]),
        .I4(\r3/t3/t0/p_1_in [0]),
        .I5(\r3/t3/t0/p_0_in [0]),
        .O(\r3/p_0_out [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[0]_i_1__2 
       (.I0(\r4/t0/t1/p_0_in [0]),
        .I1(\r4/t2/t3/p_1_in [0]),
        .I2(\r4/t1/t2/p_0_in [0]),
        .I3(k3b[0]),
        .I4(\r4/t3/t0/p_1_in [0]),
        .I5(\r4/t3/t0/p_0_in [0]),
        .O(\r4/p_0_out [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[0]_i_1__3 
       (.I0(\r5/t0/t1/p_0_in [0]),
        .I1(\r5/t2/t3/p_1_in [0]),
        .I2(\r5/t1/t2/p_0_in [0]),
        .I3(k4b[0]),
        .I4(\r5/t3/t0/p_1_in [0]),
        .I5(\r5/t3/t0/p_0_in [0]),
        .O(\r5/p_0_out [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[0]_i_1__4 
       (.I0(\r6/t0/t1/p_0_in [0]),
        .I1(\r6/t2/t3/p_1_in [0]),
        .I2(\r6/t1/t2/p_0_in [0]),
        .I3(k5b[0]),
        .I4(\r6/t3/t0/p_1_in [0]),
        .I5(\r6/t3/t0/p_0_in [0]),
        .O(\r6/p_0_out [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[0]_i_1__5 
       (.I0(\r7/t0/t1/p_0_in [0]),
        .I1(\r7/t2/t3/p_1_in [0]),
        .I2(\r7/t1/t2/p_0_in [0]),
        .I3(k6b[0]),
        .I4(\r7/t3/t0/p_1_in [0]),
        .I5(\r7/t3/t0/p_0_in [0]),
        .O(\r7/p_0_out [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[0]_i_1__6 
       (.I0(\r8/t0/t1/p_0_in [0]),
        .I1(\r8/t2/t3/p_1_in [0]),
        .I2(\r8/t1/t2/p_0_in [0]),
        .I3(k7b[0]),
        .I4(\r8/t3/t0/p_1_in [0]),
        .I5(\r8/t3/t0/p_0_in [0]),
        .O(\r8/p_0_out [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[0]_i_1__7 
       (.I0(\r9/t0/t1/p_0_in [0]),
        .I1(\r9/t2/t3/p_1_in [0]),
        .I2(\r9/t1/t2/p_0_in [0]),
        .I3(k8b[0]),
        .I4(\r9/t3/t0/p_1_in [0]),
        .I5(\r9/t3/t0/p_0_in [0]),
        .O(\r9/p_0_out [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair342" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[0]_i_1__8 
       (.I0(\a10/k3a [0]),
        .I1(\a10/k4a [0]),
        .I2(\rf/p_0_in [0]),
        .O(\rf/p_4_out [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[100]_i_1 
       (.I0(\r1/t0/t0/p_1_in [4]),
        .I1(\r1/t0/t0/p_0_in [4]),
        .I2(\r1/t2/t2/p_0_in [4]),
        .I3(\r1/t1/t1/p_0_in [4]),
        .I4(k0b[100]),
        .I5(\r1/t3/t3/p_1_in [4]),
        .O(\r1/p_0_out [100]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[100]_i_1__0 
       (.I0(\r2/t0/t0/p_1_in [4]),
        .I1(\r2/t0/t0/p_0_in [4]),
        .I2(\r2/t2/t2/p_0_in [4]),
        .I3(\r2/t1/t1/p_0_in [4]),
        .I4(k1b[100]),
        .I5(\r2/t3/t3/p_1_in [4]),
        .O(\r2/p_0_out [100]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[100]_i_1__1 
       (.I0(\r3/t0/t0/p_1_in [4]),
        .I1(\r3/t0/t0/p_0_in [4]),
        .I2(\r3/t2/t2/p_0_in [4]),
        .I3(\r3/t1/t1/p_0_in [4]),
        .I4(k2b[100]),
        .I5(\r3/t3/t3/p_1_in [4]),
        .O(\r3/p_0_out [100]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[100]_i_1__2 
       (.I0(\r4/t0/t0/p_1_in [4]),
        .I1(\r4/t0/t0/p_0_in [4]),
        .I2(\r4/t2/t2/p_0_in [4]),
        .I3(\r4/t1/t1/p_0_in [4]),
        .I4(k3b[100]),
        .I5(\r4/t3/t3/p_1_in [4]),
        .O(\r4/p_0_out [100]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[100]_i_1__3 
       (.I0(\r5/t0/t0/p_1_in [4]),
        .I1(\r5/t0/t0/p_0_in [4]),
        .I2(\r5/t2/t2/p_0_in [4]),
        .I3(\r5/t1/t1/p_0_in [4]),
        .I4(k4b[100]),
        .I5(\r5/t3/t3/p_1_in [4]),
        .O(\r5/p_0_out [100]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[100]_i_1__4 
       (.I0(\r6/t0/t0/p_1_in [4]),
        .I1(\r6/t0/t0/p_0_in [4]),
        .I2(\r6/t2/t2/p_0_in [4]),
        .I3(\r6/t1/t1/p_0_in [4]),
        .I4(k5b[100]),
        .I5(\r6/t3/t3/p_1_in [4]),
        .O(\r6/p_0_out [100]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[100]_i_1__5 
       (.I0(\r7/t0/t0/p_1_in [4]),
        .I1(\r7/t0/t0/p_0_in [4]),
        .I2(\r7/t2/t2/p_0_in [4]),
        .I3(\r7/t1/t1/p_0_in [4]),
        .I4(k6b[100]),
        .I5(\r7/t3/t3/p_1_in [4]),
        .O(\r7/p_0_out [100]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[100]_i_1__6 
       (.I0(\r8/t0/t0/p_1_in [4]),
        .I1(\r8/t0/t0/p_0_in [4]),
        .I2(\r8/t2/t2/p_0_in [4]),
        .I3(\r8/t1/t1/p_0_in [4]),
        .I4(k7b[100]),
        .I5(\r8/t3/t3/p_1_in [4]),
        .O(\r8/p_0_out [100]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[100]_i_1__7 
       (.I0(\r9/t0/t0/p_1_in [4]),
        .I1(\r9/t0/t0/p_0_in [4]),
        .I2(\r9/t2/t2/p_0_in [4]),
        .I3(\r9/t1/t1/p_0_in [4]),
        .I4(k8b[100]),
        .I5(\r9/t3/t3/p_1_in [4]),
        .O(\r9/p_0_out [100]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair338" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[100]_i_1__8 
       (.I0(\a10/k0a [4]),
        .I1(\a10/k4a [4]),
        .I2(\rf/p_3_in [4]),
        .O(\rf/p_4_out [100]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[101]_i_1 
       (.I0(\r1/t0/t0/p_1_in [5]),
        .I1(\r1/t0/t0/p_0_in [5]),
        .I2(\r1/t2/t2/p_0_in [5]),
        .I3(\r1/t1/t1/p_0_in [5]),
        .I4(k0b[101]),
        .I5(\r1/t3/t3/p_1_in [5]),
        .O(\r1/p_0_out [101]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[101]_i_1__0 
       (.I0(\r2/t0/t0/p_1_in [5]),
        .I1(\r2/t0/t0/p_0_in [5]),
        .I2(\r2/t2/t2/p_0_in [5]),
        .I3(\r2/t1/t1/p_0_in [5]),
        .I4(k1b[101]),
        .I5(\r2/t3/t3/p_1_in [5]),
        .O(\r2/p_0_out [101]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[101]_i_1__1 
       (.I0(\r3/t0/t0/p_1_in [5]),
        .I1(\r3/t0/t0/p_0_in [5]),
        .I2(\r3/t2/t2/p_0_in [5]),
        .I3(\r3/t1/t1/p_0_in [5]),
        .I4(k2b[101]),
        .I5(\r3/t3/t3/p_1_in [5]),
        .O(\r3/p_0_out [101]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[101]_i_1__2 
       (.I0(\r4/t0/t0/p_1_in [5]),
        .I1(\r4/t0/t0/p_0_in [5]),
        .I2(\r4/t2/t2/p_0_in [5]),
        .I3(\r4/t1/t1/p_0_in [5]),
        .I4(k3b[101]),
        .I5(\r4/t3/t3/p_1_in [5]),
        .O(\r4/p_0_out [101]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[101]_i_1__3 
       (.I0(\r5/t0/t0/p_1_in [5]),
        .I1(\r5/t0/t0/p_0_in [5]),
        .I2(\r5/t2/t2/p_0_in [5]),
        .I3(\r5/t1/t1/p_0_in [5]),
        .I4(k4b[101]),
        .I5(\r5/t3/t3/p_1_in [5]),
        .O(\r5/p_0_out [101]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[101]_i_1__4 
       (.I0(\r6/t0/t0/p_1_in [5]),
        .I1(\r6/t0/t0/p_0_in [5]),
        .I2(\r6/t2/t2/p_0_in [5]),
        .I3(\r6/t1/t1/p_0_in [5]),
        .I4(k5b[101]),
        .I5(\r6/t3/t3/p_1_in [5]),
        .O(\r6/p_0_out [101]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[101]_i_1__5 
       (.I0(\r7/t0/t0/p_1_in [5]),
        .I1(\r7/t0/t0/p_0_in [5]),
        .I2(\r7/t2/t2/p_0_in [5]),
        .I3(\r7/t1/t1/p_0_in [5]),
        .I4(k6b[101]),
        .I5(\r7/t3/t3/p_1_in [5]),
        .O(\r7/p_0_out [101]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[101]_i_1__6 
       (.I0(\r8/t0/t0/p_1_in [5]),
        .I1(\r8/t0/t0/p_0_in [5]),
        .I2(\r8/t2/t2/p_0_in [5]),
        .I3(\r8/t1/t1/p_0_in [5]),
        .I4(k7b[101]),
        .I5(\r8/t3/t3/p_1_in [5]),
        .O(\r8/p_0_out [101]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[101]_i_1__7 
       (.I0(\r9/t0/t0/p_1_in [5]),
        .I1(\r9/t0/t0/p_0_in [5]),
        .I2(\r9/t2/t2/p_0_in [5]),
        .I3(\r9/t1/t1/p_0_in [5]),
        .I4(k8b[101]),
        .I5(\r9/t3/t3/p_1_in [5]),
        .O(\r9/p_0_out [101]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair337" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[101]_i_1__8 
       (.I0(\a10/k0a [5]),
        .I1(\a10/k4a [5]),
        .I2(\rf/p_3_in [5]),
        .O(\rf/p_4_out [101]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[102]_i_1 
       (.I0(\r1/t0/t0/p_1_in [6]),
        .I1(\r1/t0/t0/p_0_in [6]),
        .I2(\r1/t2/t2/p_0_in [6]),
        .I3(\r1/t1/t1/p_0_in [6]),
        .I4(k0b[102]),
        .I5(\r1/t3/t3/p_1_in [6]),
        .O(\r1/p_0_out [102]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[102]_i_1__0 
       (.I0(\r2/t0/t0/p_1_in [6]),
        .I1(\r2/t0/t0/p_0_in [6]),
        .I2(\r2/t2/t2/p_0_in [6]),
        .I3(\r2/t1/t1/p_0_in [6]),
        .I4(k1b[102]),
        .I5(\r2/t3/t3/p_1_in [6]),
        .O(\r2/p_0_out [102]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[102]_i_1__1 
       (.I0(\r3/t0/t0/p_1_in [6]),
        .I1(\r3/t0/t0/p_0_in [6]),
        .I2(\r3/t2/t2/p_0_in [6]),
        .I3(\r3/t1/t1/p_0_in [6]),
        .I4(k2b[102]),
        .I5(\r3/t3/t3/p_1_in [6]),
        .O(\r3/p_0_out [102]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[102]_i_1__2 
       (.I0(\r4/t0/t0/p_1_in [6]),
        .I1(\r4/t0/t0/p_0_in [6]),
        .I2(\r4/t2/t2/p_0_in [6]),
        .I3(\r4/t1/t1/p_0_in [6]),
        .I4(k3b[102]),
        .I5(\r4/t3/t3/p_1_in [6]),
        .O(\r4/p_0_out [102]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[102]_i_1__3 
       (.I0(\r5/t0/t0/p_1_in [6]),
        .I1(\r5/t0/t0/p_0_in [6]),
        .I2(\r5/t2/t2/p_0_in [6]),
        .I3(\r5/t1/t1/p_0_in [6]),
        .I4(k4b[102]),
        .I5(\r5/t3/t3/p_1_in [6]),
        .O(\r5/p_0_out [102]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[102]_i_1__4 
       (.I0(\r6/t0/t0/p_1_in [6]),
        .I1(\r6/t0/t0/p_0_in [6]),
        .I2(\r6/t2/t2/p_0_in [6]),
        .I3(\r6/t1/t1/p_0_in [6]),
        .I4(k5b[102]),
        .I5(\r6/t3/t3/p_1_in [6]),
        .O(\r6/p_0_out [102]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[102]_i_1__5 
       (.I0(\r7/t0/t0/p_1_in [6]),
        .I1(\r7/t0/t0/p_0_in [6]),
        .I2(\r7/t2/t2/p_0_in [6]),
        .I3(\r7/t1/t1/p_0_in [6]),
        .I4(k6b[102]),
        .I5(\r7/t3/t3/p_1_in [6]),
        .O(\r7/p_0_out [102]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[102]_i_1__6 
       (.I0(\r8/t0/t0/p_1_in [6]),
        .I1(\r8/t0/t0/p_0_in [6]),
        .I2(\r8/t2/t2/p_0_in [6]),
        .I3(\r8/t1/t1/p_0_in [6]),
        .I4(k7b[102]),
        .I5(\r8/t3/t3/p_1_in [6]),
        .O(\r8/p_0_out [102]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[102]_i_1__7 
       (.I0(\r9/t0/t0/p_1_in [6]),
        .I1(\r9/t0/t0/p_0_in [6]),
        .I2(\r9/t2/t2/p_0_in [6]),
        .I3(\r9/t1/t1/p_0_in [6]),
        .I4(k8b[102]),
        .I5(\r9/t3/t3/p_1_in [6]),
        .O(\r9/p_0_out [102]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair336" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[102]_i_1__8 
       (.I0(\a10/k0a [6]),
        .I1(\a10/k4a [6]),
        .I2(\rf/p_3_in [6]),
        .O(\rf/p_4_out [102]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[103]_i_1 
       (.I0(\r1/t0/t0/p_1_in [7]),
        .I1(\r1/t0/t0/p_0_in [7]),
        .I2(\r1/t2/t2/p_0_in [7]),
        .I3(\r1/t1/t1/p_0_in [7]),
        .I4(k0b[103]),
        .I5(\r1/t3/t3/p_1_in [7]),
        .O(\r1/p_0_out [103]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[103]_i_1__0 
       (.I0(\r2/t0/t0/p_1_in [7]),
        .I1(\r2/t0/t0/p_0_in [7]),
        .I2(\r2/t2/t2/p_0_in [7]),
        .I3(\r2/t1/t1/p_0_in [7]),
        .I4(k1b[103]),
        .I5(\r2/t3/t3/p_1_in [7]),
        .O(\r2/p_0_out [103]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[103]_i_1__1 
       (.I0(\r3/t0/t0/p_1_in [7]),
        .I1(\r3/t0/t0/p_0_in [7]),
        .I2(\r3/t2/t2/p_0_in [7]),
        .I3(\r3/t1/t1/p_0_in [7]),
        .I4(k2b[103]),
        .I5(\r3/t3/t3/p_1_in [7]),
        .O(\r3/p_0_out [103]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[103]_i_1__2 
       (.I0(\r4/t0/t0/p_1_in [7]),
        .I1(\r4/t0/t0/p_0_in [7]),
        .I2(\r4/t2/t2/p_0_in [7]),
        .I3(\r4/t1/t1/p_0_in [7]),
        .I4(k3b[103]),
        .I5(\r4/t3/t3/p_1_in [7]),
        .O(\r4/p_0_out [103]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[103]_i_1__3 
       (.I0(\r5/t0/t0/p_1_in [7]),
        .I1(\r5/t0/t0/p_0_in [7]),
        .I2(\r5/t2/t2/p_0_in [7]),
        .I3(\r5/t1/t1/p_0_in [7]),
        .I4(k4b[103]),
        .I5(\r5/t3/t3/p_1_in [7]),
        .O(\r5/p_0_out [103]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[103]_i_1__4 
       (.I0(\r6/t0/t0/p_1_in [7]),
        .I1(\r6/t0/t0/p_0_in [7]),
        .I2(\r6/t2/t2/p_0_in [7]),
        .I3(\r6/t1/t1/p_0_in [7]),
        .I4(k5b[103]),
        .I5(\r6/t3/t3/p_1_in [7]),
        .O(\r6/p_0_out [103]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[103]_i_1__5 
       (.I0(\r7/t0/t0/p_1_in [7]),
        .I1(\r7/t0/t0/p_0_in [7]),
        .I2(\r7/t2/t2/p_0_in [7]),
        .I3(\r7/t1/t1/p_0_in [7]),
        .I4(k6b[103]),
        .I5(\r7/t3/t3/p_1_in [7]),
        .O(\r7/p_0_out [103]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[103]_i_1__6 
       (.I0(\r8/t0/t0/p_1_in [7]),
        .I1(\r8/t0/t0/p_0_in [7]),
        .I2(\r8/t2/t2/p_0_in [7]),
        .I3(\r8/t1/t1/p_0_in [7]),
        .I4(k7b[103]),
        .I5(\r8/t3/t3/p_1_in [7]),
        .O(\r8/p_0_out [103]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[103]_i_1__7 
       (.I0(\r9/t0/t0/p_1_in [7]),
        .I1(\r9/t0/t0/p_0_in [7]),
        .I2(\r9/t2/t2/p_0_in [7]),
        .I3(\r9/t1/t1/p_0_in [7]),
        .I4(k8b[103]),
        .I5(\r9/t3/t3/p_1_in [7]),
        .O(\r9/p_0_out [103]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair335" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[103]_i_1__8 
       (.I0(\a10/k0a [7]),
        .I1(\a10/k4a [7]),
        .I2(\rf/p_3_in [7]),
        .O(\rf/p_4_out [103]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[104]_i_1 
       (.I0(\r1/t0/t0/p_0_in [0]),
        .I1(\r1/t2/t2/p_1_in [0]),
        .I2(\r1/t1/t1/p_0_in [0]),
        .I3(k0b[104]),
        .I4(\r1/t3/t3/p_1_in [0]),
        .I5(\r1/t3/t3/p_0_in [0]),
        .O(\r1/p_0_out [104]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[104]_i_1__0 
       (.I0(\r2/t0/t0/p_0_in [0]),
        .I1(\r2/t2/t2/p_1_in [0]),
        .I2(\r2/t1/t1/p_0_in [0]),
        .I3(k1b[104]),
        .I4(\r2/t3/t3/p_1_in [0]),
        .I5(\r2/t3/t3/p_0_in [0]),
        .O(\r2/p_0_out [104]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[104]_i_1__1 
       (.I0(\r3/t0/t0/p_0_in [0]),
        .I1(\r3/t2/t2/p_1_in [0]),
        .I2(\r3/t1/t1/p_0_in [0]),
        .I3(k2b[104]),
        .I4(\r3/t3/t3/p_1_in [0]),
        .I5(\r3/t3/t3/p_0_in [0]),
        .O(\r3/p_0_out [104]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[104]_i_1__2 
       (.I0(\r4/t0/t0/p_0_in [0]),
        .I1(\r4/t2/t2/p_1_in [0]),
        .I2(\r4/t1/t1/p_0_in [0]),
        .I3(k3b[104]),
        .I4(\r4/t3/t3/p_1_in [0]),
        .I5(\r4/t3/t3/p_0_in [0]),
        .O(\r4/p_0_out [104]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[104]_i_1__3 
       (.I0(\r5/t0/t0/p_0_in [0]),
        .I1(\r5/t2/t2/p_1_in [0]),
        .I2(\r5/t1/t1/p_0_in [0]),
        .I3(k4b[104]),
        .I4(\r5/t3/t3/p_1_in [0]),
        .I5(\r5/t3/t3/p_0_in [0]),
        .O(\r5/p_0_out [104]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[104]_i_1__4 
       (.I0(\r6/t0/t0/p_0_in [0]),
        .I1(\r6/t2/t2/p_1_in [0]),
        .I2(\r6/t1/t1/p_0_in [0]),
        .I3(k5b[104]),
        .I4(\r6/t3/t3/p_1_in [0]),
        .I5(\r6/t3/t3/p_0_in [0]),
        .O(\r6/p_0_out [104]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[104]_i_1__5 
       (.I0(\r7/t0/t0/p_0_in [0]),
        .I1(\r7/t2/t2/p_1_in [0]),
        .I2(\r7/t1/t1/p_0_in [0]),
        .I3(k6b[104]),
        .I4(\r7/t3/t3/p_1_in [0]),
        .I5(\r7/t3/t3/p_0_in [0]),
        .O(\r7/p_0_out [104]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[104]_i_1__6 
       (.I0(\r8/t0/t0/p_0_in [0]),
        .I1(\r8/t2/t2/p_1_in [0]),
        .I2(\r8/t1/t1/p_0_in [0]),
        .I3(k7b[104]),
        .I4(\r8/t3/t3/p_1_in [0]),
        .I5(\r8/t3/t3/p_0_in [0]),
        .O(\r8/p_0_out [104]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[104]_i_1__7 
       (.I0(\r9/t0/t0/p_0_in [0]),
        .I1(\r9/t2/t2/p_1_in [0]),
        .I2(\r9/t1/t1/p_0_in [0]),
        .I3(k8b[104]),
        .I4(\r9/t3/t3/p_1_in [0]),
        .I5(\r9/t3/t3/p_0_in [0]),
        .O(\r9/p_0_out [104]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair334" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[104]_i_1__8 
       (.I0(\a10/k0a [8]),
        .I1(\a10/k4a [8]),
        .I2(\rf/p_3_in [8]),
        .O(\rf/p_4_out [104]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[105]_i_1 
       (.I0(\r1/t0/t0/p_0_in [1]),
        .I1(\r1/t2/t2/p_1_in [1]),
        .I2(\r1/t1/t1/p_0_in [1]),
        .I3(k0b[105]),
        .I4(\r1/t3/t3/p_1_in [1]),
        .I5(\r1/t3/t3/p_0_in [1]),
        .O(\r1/p_0_out [105]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[105]_i_1__0 
       (.I0(\r2/t0/t0/p_0_in [1]),
        .I1(\r2/t2/t2/p_1_in [1]),
        .I2(\r2/t1/t1/p_0_in [1]),
        .I3(k1b[105]),
        .I4(\r2/t3/t3/p_1_in [1]),
        .I5(\r2/t3/t3/p_0_in [1]),
        .O(\r2/p_0_out [105]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[105]_i_1__1 
       (.I0(\r3/t0/t0/p_0_in [1]),
        .I1(\r3/t2/t2/p_1_in [1]),
        .I2(\r3/t1/t1/p_0_in [1]),
        .I3(k2b[105]),
        .I4(\r3/t3/t3/p_1_in [1]),
        .I5(\r3/t3/t3/p_0_in [1]),
        .O(\r3/p_0_out [105]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[105]_i_1__2 
       (.I0(\r4/t0/t0/p_0_in [1]),
        .I1(\r4/t2/t2/p_1_in [1]),
        .I2(\r4/t1/t1/p_0_in [1]),
        .I3(k3b[105]),
        .I4(\r4/t3/t3/p_1_in [1]),
        .I5(\r4/t3/t3/p_0_in [1]),
        .O(\r4/p_0_out [105]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[105]_i_1__3 
       (.I0(\r5/t0/t0/p_0_in [1]),
        .I1(\r5/t2/t2/p_1_in [1]),
        .I2(\r5/t1/t1/p_0_in [1]),
        .I3(k4b[105]),
        .I4(\r5/t3/t3/p_1_in [1]),
        .I5(\r5/t3/t3/p_0_in [1]),
        .O(\r5/p_0_out [105]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[105]_i_1__4 
       (.I0(\r6/t0/t0/p_0_in [1]),
        .I1(\r6/t2/t2/p_1_in [1]),
        .I2(\r6/t1/t1/p_0_in [1]),
        .I3(k5b[105]),
        .I4(\r6/t3/t3/p_1_in [1]),
        .I5(\r6/t3/t3/p_0_in [1]),
        .O(\r6/p_0_out [105]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[105]_i_1__5 
       (.I0(\r7/t0/t0/p_0_in [1]),
        .I1(\r7/t2/t2/p_1_in [1]),
        .I2(\r7/t1/t1/p_0_in [1]),
        .I3(k6b[105]),
        .I4(\r7/t3/t3/p_1_in [1]),
        .I5(\r7/t3/t3/p_0_in [1]),
        .O(\r7/p_0_out [105]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[105]_i_1__6 
       (.I0(\r8/t0/t0/p_0_in [1]),
        .I1(\r8/t2/t2/p_1_in [1]),
        .I2(\r8/t1/t1/p_0_in [1]),
        .I3(k7b[105]),
        .I4(\r8/t3/t3/p_1_in [1]),
        .I5(\r8/t3/t3/p_0_in [1]),
        .O(\r8/p_0_out [105]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[105]_i_1__7 
       (.I0(\r9/t0/t0/p_0_in [1]),
        .I1(\r9/t2/t2/p_1_in [1]),
        .I2(\r9/t1/t1/p_0_in [1]),
        .I3(k8b[105]),
        .I4(\r9/t3/t3/p_1_in [1]),
        .I5(\r9/t3/t3/p_0_in [1]),
        .O(\r9/p_0_out [105]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair333" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[105]_i_1__8 
       (.I0(\a10/k0a [9]),
        .I1(\a10/k4a [9]),
        .I2(\rf/p_3_in [9]),
        .O(\rf/p_4_out [105]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[106]_i_1 
       (.I0(\r1/t0/t0/p_0_in [2]),
        .I1(\r1/t2/t2/p_1_in [2]),
        .I2(\r1/t1/t1/p_0_in [2]),
        .I3(k0b[106]),
        .I4(\r1/t3/t3/p_1_in [2]),
        .I5(\r1/t3/t3/p_0_in [2]),
        .O(\r1/p_0_out [106]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[106]_i_1__0 
       (.I0(\r2/t0/t0/p_0_in [2]),
        .I1(\r2/t2/t2/p_1_in [2]),
        .I2(\r2/t1/t1/p_0_in [2]),
        .I3(k1b[106]),
        .I4(\r2/t3/t3/p_1_in [2]),
        .I5(\r2/t3/t3/p_0_in [2]),
        .O(\r2/p_0_out [106]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[106]_i_1__1 
       (.I0(\r3/t0/t0/p_0_in [2]),
        .I1(\r3/t2/t2/p_1_in [2]),
        .I2(\r3/t1/t1/p_0_in [2]),
        .I3(k2b[106]),
        .I4(\r3/t3/t3/p_1_in [2]),
        .I5(\r3/t3/t3/p_0_in [2]),
        .O(\r3/p_0_out [106]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[106]_i_1__2 
       (.I0(\r4/t0/t0/p_0_in [2]),
        .I1(\r4/t2/t2/p_1_in [2]),
        .I2(\r4/t1/t1/p_0_in [2]),
        .I3(k3b[106]),
        .I4(\r4/t3/t3/p_1_in [2]),
        .I5(\r4/t3/t3/p_0_in [2]),
        .O(\r4/p_0_out [106]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[106]_i_1__3 
       (.I0(\r5/t0/t0/p_0_in [2]),
        .I1(\r5/t2/t2/p_1_in [2]),
        .I2(\r5/t1/t1/p_0_in [2]),
        .I3(k4b[106]),
        .I4(\r5/t3/t3/p_1_in [2]),
        .I5(\r5/t3/t3/p_0_in [2]),
        .O(\r5/p_0_out [106]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[106]_i_1__4 
       (.I0(\r6/t0/t0/p_0_in [2]),
        .I1(\r6/t2/t2/p_1_in [2]),
        .I2(\r6/t1/t1/p_0_in [2]),
        .I3(k5b[106]),
        .I4(\r6/t3/t3/p_1_in [2]),
        .I5(\r6/t3/t3/p_0_in [2]),
        .O(\r6/p_0_out [106]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[106]_i_1__5 
       (.I0(\r7/t0/t0/p_0_in [2]),
        .I1(\r7/t2/t2/p_1_in [2]),
        .I2(\r7/t1/t1/p_0_in [2]),
        .I3(k6b[106]),
        .I4(\r7/t3/t3/p_1_in [2]),
        .I5(\r7/t3/t3/p_0_in [2]),
        .O(\r7/p_0_out [106]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[106]_i_1__6 
       (.I0(\r8/t0/t0/p_0_in [2]),
        .I1(\r8/t2/t2/p_1_in [2]),
        .I2(\r8/t1/t1/p_0_in [2]),
        .I3(k7b[106]),
        .I4(\r8/t3/t3/p_1_in [2]),
        .I5(\r8/t3/t3/p_0_in [2]),
        .O(\r8/p_0_out [106]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[106]_i_1__7 
       (.I0(\r9/t0/t0/p_0_in [2]),
        .I1(\r9/t2/t2/p_1_in [2]),
        .I2(\r9/t1/t1/p_0_in [2]),
        .I3(k8b[106]),
        .I4(\r9/t3/t3/p_1_in [2]),
        .I5(\r9/t3/t3/p_0_in [2]),
        .O(\r9/p_0_out [106]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair332" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[106]_i_1__8 
       (.I0(\a10/k0a [10]),
        .I1(\a10/k4a [10]),
        .I2(\rf/p_3_in [10]),
        .O(\rf/p_4_out [106]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[107]_i_1 
       (.I0(\r1/t0/t0/p_0_in [3]),
        .I1(\r1/t2/t2/p_1_in [3]),
        .I2(\r1/t1/t1/p_0_in [3]),
        .I3(k0b[107]),
        .I4(\r1/t3/t3/p_1_in [3]),
        .I5(\r1/t3/t3/p_0_in [3]),
        .O(\r1/p_0_out [107]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[107]_i_1__0 
       (.I0(\r2/t0/t0/p_0_in [3]),
        .I1(\r2/t2/t2/p_1_in [3]),
        .I2(\r2/t1/t1/p_0_in [3]),
        .I3(k1b[107]),
        .I4(\r2/t3/t3/p_1_in [3]),
        .I5(\r2/t3/t3/p_0_in [3]),
        .O(\r2/p_0_out [107]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[107]_i_1__1 
       (.I0(\r3/t0/t0/p_0_in [3]),
        .I1(\r3/t2/t2/p_1_in [3]),
        .I2(\r3/t1/t1/p_0_in [3]),
        .I3(k2b[107]),
        .I4(\r3/t3/t3/p_1_in [3]),
        .I5(\r3/t3/t3/p_0_in [3]),
        .O(\r3/p_0_out [107]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[107]_i_1__2 
       (.I0(\r4/t0/t0/p_0_in [3]),
        .I1(\r4/t2/t2/p_1_in [3]),
        .I2(\r4/t1/t1/p_0_in [3]),
        .I3(k3b[107]),
        .I4(\r4/t3/t3/p_1_in [3]),
        .I5(\r4/t3/t3/p_0_in [3]),
        .O(\r4/p_0_out [107]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[107]_i_1__3 
       (.I0(\r5/t0/t0/p_0_in [3]),
        .I1(\r5/t2/t2/p_1_in [3]),
        .I2(\r5/t1/t1/p_0_in [3]),
        .I3(k4b[107]),
        .I4(\r5/t3/t3/p_1_in [3]),
        .I5(\r5/t3/t3/p_0_in [3]),
        .O(\r5/p_0_out [107]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[107]_i_1__4 
       (.I0(\r6/t0/t0/p_0_in [3]),
        .I1(\r6/t2/t2/p_1_in [3]),
        .I2(\r6/t1/t1/p_0_in [3]),
        .I3(k5b[107]),
        .I4(\r6/t3/t3/p_1_in [3]),
        .I5(\r6/t3/t3/p_0_in [3]),
        .O(\r6/p_0_out [107]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[107]_i_1__5 
       (.I0(\r7/t0/t0/p_0_in [3]),
        .I1(\r7/t2/t2/p_1_in [3]),
        .I2(\r7/t1/t1/p_0_in [3]),
        .I3(k6b[107]),
        .I4(\r7/t3/t3/p_1_in [3]),
        .I5(\r7/t3/t3/p_0_in [3]),
        .O(\r7/p_0_out [107]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[107]_i_1__6 
       (.I0(\r8/t0/t0/p_0_in [3]),
        .I1(\r8/t2/t2/p_1_in [3]),
        .I2(\r8/t1/t1/p_0_in [3]),
        .I3(k7b[107]),
        .I4(\r8/t3/t3/p_1_in [3]),
        .I5(\r8/t3/t3/p_0_in [3]),
        .O(\r8/p_0_out [107]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[107]_i_1__7 
       (.I0(\r9/t0/t0/p_0_in [3]),
        .I1(\r9/t2/t2/p_1_in [3]),
        .I2(\r9/t1/t1/p_0_in [3]),
        .I3(k8b[107]),
        .I4(\r9/t3/t3/p_1_in [3]),
        .I5(\r9/t3/t3/p_0_in [3]),
        .O(\r9/p_0_out [107]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair331" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[107]_i_1__8 
       (.I0(\a10/k0a [11]),
        .I1(\a10/k4a [11]),
        .I2(\rf/p_3_in [11]),
        .O(\rf/p_4_out [107]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[108]_i_1 
       (.I0(\r1/t0/t0/p_0_in [4]),
        .I1(\r1/t2/t2/p_1_in [4]),
        .I2(\r1/t1/t1/p_0_in [4]),
        .I3(k0b[108]),
        .I4(\r1/t3/t3/p_1_in [4]),
        .I5(\r1/t3/t3/p_0_in [4]),
        .O(\r1/p_0_out [108]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[108]_i_1__0 
       (.I0(\r2/t0/t0/p_0_in [4]),
        .I1(\r2/t2/t2/p_1_in [4]),
        .I2(\r2/t1/t1/p_0_in [4]),
        .I3(k1b[108]),
        .I4(\r2/t3/t3/p_1_in [4]),
        .I5(\r2/t3/t3/p_0_in [4]),
        .O(\r2/p_0_out [108]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[108]_i_1__1 
       (.I0(\r3/t0/t0/p_0_in [4]),
        .I1(\r3/t2/t2/p_1_in [4]),
        .I2(\r3/t1/t1/p_0_in [4]),
        .I3(k2b[108]),
        .I4(\r3/t3/t3/p_1_in [4]),
        .I5(\r3/t3/t3/p_0_in [4]),
        .O(\r3/p_0_out [108]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[108]_i_1__2 
       (.I0(\r4/t0/t0/p_0_in [4]),
        .I1(\r4/t2/t2/p_1_in [4]),
        .I2(\r4/t1/t1/p_0_in [4]),
        .I3(k3b[108]),
        .I4(\r4/t3/t3/p_1_in [4]),
        .I5(\r4/t3/t3/p_0_in [4]),
        .O(\r4/p_0_out [108]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[108]_i_1__3 
       (.I0(\r5/t0/t0/p_0_in [4]),
        .I1(\r5/t2/t2/p_1_in [4]),
        .I2(\r5/t1/t1/p_0_in [4]),
        .I3(k4b[108]),
        .I4(\r5/t3/t3/p_1_in [4]),
        .I5(\r5/t3/t3/p_0_in [4]),
        .O(\r5/p_0_out [108]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[108]_i_1__4 
       (.I0(\r6/t0/t0/p_0_in [4]),
        .I1(\r6/t2/t2/p_1_in [4]),
        .I2(\r6/t1/t1/p_0_in [4]),
        .I3(k5b[108]),
        .I4(\r6/t3/t3/p_1_in [4]),
        .I5(\r6/t3/t3/p_0_in [4]),
        .O(\r6/p_0_out [108]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[108]_i_1__5 
       (.I0(\r7/t0/t0/p_0_in [4]),
        .I1(\r7/t2/t2/p_1_in [4]),
        .I2(\r7/t1/t1/p_0_in [4]),
        .I3(k6b[108]),
        .I4(\r7/t3/t3/p_1_in [4]),
        .I5(\r7/t3/t3/p_0_in [4]),
        .O(\r7/p_0_out [108]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[108]_i_1__6 
       (.I0(\r8/t0/t0/p_0_in [4]),
        .I1(\r8/t2/t2/p_1_in [4]),
        .I2(\r8/t1/t1/p_0_in [4]),
        .I3(k7b[108]),
        .I4(\r8/t3/t3/p_1_in [4]),
        .I5(\r8/t3/t3/p_0_in [4]),
        .O(\r8/p_0_out [108]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[108]_i_1__7 
       (.I0(\r9/t0/t0/p_0_in [4]),
        .I1(\r9/t2/t2/p_1_in [4]),
        .I2(\r9/t1/t1/p_0_in [4]),
        .I3(k8b[108]),
        .I4(\r9/t3/t3/p_1_in [4]),
        .I5(\r9/t3/t3/p_0_in [4]),
        .O(\r9/p_0_out [108]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair330" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[108]_i_1__8 
       (.I0(\a10/k0a [12]),
        .I1(\a10/k4a [12]),
        .I2(\rf/p_3_in [12]),
        .O(\rf/p_4_out [108]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[109]_i_1 
       (.I0(\r1/t0/t0/p_0_in [5]),
        .I1(\r1/t2/t2/p_1_in [5]),
        .I2(\r1/t1/t1/p_0_in [5]),
        .I3(k0b[109]),
        .I4(\r1/t3/t3/p_1_in [5]),
        .I5(\r1/t3/t3/p_0_in [5]),
        .O(\r1/p_0_out [109]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[109]_i_1__0 
       (.I0(\r2/t0/t0/p_0_in [5]),
        .I1(\r2/t2/t2/p_1_in [5]),
        .I2(\r2/t1/t1/p_0_in [5]),
        .I3(k1b[109]),
        .I4(\r2/t3/t3/p_1_in [5]),
        .I5(\r2/t3/t3/p_0_in [5]),
        .O(\r2/p_0_out [109]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[109]_i_1__1 
       (.I0(\r3/t0/t0/p_0_in [5]),
        .I1(\r3/t2/t2/p_1_in [5]),
        .I2(\r3/t1/t1/p_0_in [5]),
        .I3(k2b[109]),
        .I4(\r3/t3/t3/p_1_in [5]),
        .I5(\r3/t3/t3/p_0_in [5]),
        .O(\r3/p_0_out [109]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[109]_i_1__2 
       (.I0(\r4/t0/t0/p_0_in [5]),
        .I1(\r4/t2/t2/p_1_in [5]),
        .I2(\r4/t1/t1/p_0_in [5]),
        .I3(k3b[109]),
        .I4(\r4/t3/t3/p_1_in [5]),
        .I5(\r4/t3/t3/p_0_in [5]),
        .O(\r4/p_0_out [109]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[109]_i_1__3 
       (.I0(\r5/t0/t0/p_0_in [5]),
        .I1(\r5/t2/t2/p_1_in [5]),
        .I2(\r5/t1/t1/p_0_in [5]),
        .I3(k4b[109]),
        .I4(\r5/t3/t3/p_1_in [5]),
        .I5(\r5/t3/t3/p_0_in [5]),
        .O(\r5/p_0_out [109]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[109]_i_1__4 
       (.I0(\r6/t0/t0/p_0_in [5]),
        .I1(\r6/t2/t2/p_1_in [5]),
        .I2(\r6/t1/t1/p_0_in [5]),
        .I3(k5b[109]),
        .I4(\r6/t3/t3/p_1_in [5]),
        .I5(\r6/t3/t3/p_0_in [5]),
        .O(\r6/p_0_out [109]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[109]_i_1__5 
       (.I0(\r7/t0/t0/p_0_in [5]),
        .I1(\r7/t2/t2/p_1_in [5]),
        .I2(\r7/t1/t1/p_0_in [5]),
        .I3(k6b[109]),
        .I4(\r7/t3/t3/p_1_in [5]),
        .I5(\r7/t3/t3/p_0_in [5]),
        .O(\r7/p_0_out [109]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[109]_i_1__6 
       (.I0(\r8/t0/t0/p_0_in [5]),
        .I1(\r8/t2/t2/p_1_in [5]),
        .I2(\r8/t1/t1/p_0_in [5]),
        .I3(k7b[109]),
        .I4(\r8/t3/t3/p_1_in [5]),
        .I5(\r8/t3/t3/p_0_in [5]),
        .O(\r8/p_0_out [109]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[109]_i_1__7 
       (.I0(\r9/t0/t0/p_0_in [5]),
        .I1(\r9/t2/t2/p_1_in [5]),
        .I2(\r9/t1/t1/p_0_in [5]),
        .I3(k8b[109]),
        .I4(\r9/t3/t3/p_1_in [5]),
        .I5(\r9/t3/t3/p_0_in [5]),
        .O(\r9/p_0_out [109]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair329" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[109]_i_1__8 
       (.I0(\a10/k0a [13]),
        .I1(\a10/k4a [13]),
        .I2(\rf/p_3_in [13]),
        .O(\rf/p_4_out [109]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[10]_i_1 
       (.I0(\r1/t0/t1/p_0_in [2]),
        .I1(\r1/t2/t3/p_1_in [2]),
        .I2(\r1/t2/t3/p_0_in [2]),
        .I3(\r1/t1/t2/p_1_in [2]),
        .I4(k0b[10]),
        .I5(\r1/t3/t0/p_0_in [2]),
        .O(\r1/p_0_out [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[10]_i_1__0 
       (.I0(\r2/t0/t1/p_0_in [2]),
        .I1(\r2/t2/t3/p_1_in [2]),
        .I2(\r2/t2/t3/p_0_in [2]),
        .I3(\r2/t1/t2/p_1_in [2]),
        .I4(k1b[10]),
        .I5(\r2/t3/t0/p_0_in [2]),
        .O(\r2/p_0_out [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[10]_i_1__1 
       (.I0(\r3/t0/t1/p_0_in [2]),
        .I1(\r3/t2/t3/p_1_in [2]),
        .I2(\r3/t2/t3/p_0_in [2]),
        .I3(\r3/t1/t2/p_1_in [2]),
        .I4(k2b[10]),
        .I5(\r3/t3/t0/p_0_in [2]),
        .O(\r3/p_0_out [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[10]_i_1__2 
       (.I0(\r4/t0/t1/p_0_in [2]),
        .I1(\r4/t2/t3/p_1_in [2]),
        .I2(\r4/t2/t3/p_0_in [2]),
        .I3(\r4/t1/t2/p_1_in [2]),
        .I4(k3b[10]),
        .I5(\r4/t3/t0/p_0_in [2]),
        .O(\r4/p_0_out [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[10]_i_1__3 
       (.I0(\r5/t0/t1/p_0_in [2]),
        .I1(\r5/t2/t3/p_1_in [2]),
        .I2(\r5/t2/t3/p_0_in [2]),
        .I3(\r5/t1/t2/p_1_in [2]),
        .I4(k4b[10]),
        .I5(\r5/t3/t0/p_0_in [2]),
        .O(\r5/p_0_out [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[10]_i_1__4 
       (.I0(\r6/t0/t1/p_0_in [2]),
        .I1(\r6/t2/t3/p_1_in [2]),
        .I2(\r6/t2/t3/p_0_in [2]),
        .I3(\r6/t1/t2/p_1_in [2]),
        .I4(k5b[10]),
        .I5(\r6/t3/t0/p_0_in [2]),
        .O(\r6/p_0_out [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[10]_i_1__5 
       (.I0(\r7/t0/t1/p_0_in [2]),
        .I1(\r7/t2/t3/p_1_in [2]),
        .I2(\r7/t2/t3/p_0_in [2]),
        .I3(\r7/t1/t2/p_1_in [2]),
        .I4(k6b[10]),
        .I5(\r7/t3/t0/p_0_in [2]),
        .O(\r7/p_0_out [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[10]_i_1__6 
       (.I0(\r8/t0/t1/p_0_in [2]),
        .I1(\r8/t2/t3/p_1_in [2]),
        .I2(\r8/t2/t3/p_0_in [2]),
        .I3(\r8/t1/t2/p_1_in [2]),
        .I4(k7b[10]),
        .I5(\r8/t3/t0/p_0_in [2]),
        .O(\r8/p_0_out [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[10]_i_1__7 
       (.I0(\r9/t0/t1/p_0_in [2]),
        .I1(\r9/t2/t3/p_1_in [2]),
        .I2(\r9/t2/t3/p_0_in [2]),
        .I3(\r9/t1/t2/p_1_in [2]),
        .I4(k8b[10]),
        .I5(\r9/t3/t0/p_0_in [2]),
        .O(\r9/p_0_out [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair332" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[10]_i_1__8 
       (.I0(\a10/k3a [10]),
        .I1(\a10/k4a [10]),
        .I2(\rf/p_0_in [10]),
        .O(\rf/p_4_out [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[110]_i_1 
       (.I0(\r1/t0/t0/p_0_in [6]),
        .I1(\r1/t2/t2/p_1_in [6]),
        .I2(\r1/t1/t1/p_0_in [6]),
        .I3(k0b[110]),
        .I4(\r1/t3/t3/p_1_in [6]),
        .I5(\r1/t3/t3/p_0_in [6]),
        .O(\r1/p_0_out [110]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[110]_i_1__0 
       (.I0(\r2/t0/t0/p_0_in [6]),
        .I1(\r2/t2/t2/p_1_in [6]),
        .I2(\r2/t1/t1/p_0_in [6]),
        .I3(k1b[110]),
        .I4(\r2/t3/t3/p_1_in [6]),
        .I5(\r2/t3/t3/p_0_in [6]),
        .O(\r2/p_0_out [110]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[110]_i_1__1 
       (.I0(\r3/t0/t0/p_0_in [6]),
        .I1(\r3/t2/t2/p_1_in [6]),
        .I2(\r3/t1/t1/p_0_in [6]),
        .I3(k2b[110]),
        .I4(\r3/t3/t3/p_1_in [6]),
        .I5(\r3/t3/t3/p_0_in [6]),
        .O(\r3/p_0_out [110]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[110]_i_1__2 
       (.I0(\r4/t0/t0/p_0_in [6]),
        .I1(\r4/t2/t2/p_1_in [6]),
        .I2(\r4/t1/t1/p_0_in [6]),
        .I3(k3b[110]),
        .I4(\r4/t3/t3/p_1_in [6]),
        .I5(\r4/t3/t3/p_0_in [6]),
        .O(\r4/p_0_out [110]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[110]_i_1__3 
       (.I0(\r5/t0/t0/p_0_in [6]),
        .I1(\r5/t2/t2/p_1_in [6]),
        .I2(\r5/t1/t1/p_0_in [6]),
        .I3(k4b[110]),
        .I4(\r5/t3/t3/p_1_in [6]),
        .I5(\r5/t3/t3/p_0_in [6]),
        .O(\r5/p_0_out [110]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[110]_i_1__4 
       (.I0(\r6/t0/t0/p_0_in [6]),
        .I1(\r6/t2/t2/p_1_in [6]),
        .I2(\r6/t1/t1/p_0_in [6]),
        .I3(k5b[110]),
        .I4(\r6/t3/t3/p_1_in [6]),
        .I5(\r6/t3/t3/p_0_in [6]),
        .O(\r6/p_0_out [110]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[110]_i_1__5 
       (.I0(\r7/t0/t0/p_0_in [6]),
        .I1(\r7/t2/t2/p_1_in [6]),
        .I2(\r7/t1/t1/p_0_in [6]),
        .I3(k6b[110]),
        .I4(\r7/t3/t3/p_1_in [6]),
        .I5(\r7/t3/t3/p_0_in [6]),
        .O(\r7/p_0_out [110]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[110]_i_1__6 
       (.I0(\r8/t0/t0/p_0_in [6]),
        .I1(\r8/t2/t2/p_1_in [6]),
        .I2(\r8/t1/t1/p_0_in [6]),
        .I3(k7b[110]),
        .I4(\r8/t3/t3/p_1_in [6]),
        .I5(\r8/t3/t3/p_0_in [6]),
        .O(\r8/p_0_out [110]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[110]_i_1__7 
       (.I0(\r9/t0/t0/p_0_in [6]),
        .I1(\r9/t2/t2/p_1_in [6]),
        .I2(\r9/t1/t1/p_0_in [6]),
        .I3(k8b[110]),
        .I4(\r9/t3/t3/p_1_in [6]),
        .I5(\r9/t3/t3/p_0_in [6]),
        .O(\r9/p_0_out [110]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair328" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[110]_i_1__8 
       (.I0(\a10/k0a [14]),
        .I1(\a10/k4a [14]),
        .I2(\rf/p_3_in [14]),
        .O(\rf/p_4_out [110]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[111]_i_1 
       (.I0(\r1/t0/t0/p_0_in [7]),
        .I1(\r1/t2/t2/p_1_in [7]),
        .I2(\r1/t1/t1/p_0_in [7]),
        .I3(k0b[111]),
        .I4(\r1/t3/t3/p_1_in [7]),
        .I5(\r1/t3/t3/p_0_in [7]),
        .O(\r1/p_0_out [111]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[111]_i_1__0 
       (.I0(\r2/t0/t0/p_0_in [7]),
        .I1(\r2/t2/t2/p_1_in [7]),
        .I2(\r2/t1/t1/p_0_in [7]),
        .I3(k1b[111]),
        .I4(\r2/t3/t3/p_1_in [7]),
        .I5(\r2/t3/t3/p_0_in [7]),
        .O(\r2/p_0_out [111]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[111]_i_1__1 
       (.I0(\r3/t0/t0/p_0_in [7]),
        .I1(\r3/t2/t2/p_1_in [7]),
        .I2(\r3/t1/t1/p_0_in [7]),
        .I3(k2b[111]),
        .I4(\r3/t3/t3/p_1_in [7]),
        .I5(\r3/t3/t3/p_0_in [7]),
        .O(\r3/p_0_out [111]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[111]_i_1__2 
       (.I0(\r4/t0/t0/p_0_in [7]),
        .I1(\r4/t2/t2/p_1_in [7]),
        .I2(\r4/t1/t1/p_0_in [7]),
        .I3(k3b[111]),
        .I4(\r4/t3/t3/p_1_in [7]),
        .I5(\r4/t3/t3/p_0_in [7]),
        .O(\r4/p_0_out [111]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[111]_i_1__3 
       (.I0(\r5/t0/t0/p_0_in [7]),
        .I1(\r5/t2/t2/p_1_in [7]),
        .I2(\r5/t1/t1/p_0_in [7]),
        .I3(k4b[111]),
        .I4(\r5/t3/t3/p_1_in [7]),
        .I5(\r5/t3/t3/p_0_in [7]),
        .O(\r5/p_0_out [111]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[111]_i_1__4 
       (.I0(\r6/t0/t0/p_0_in [7]),
        .I1(\r6/t2/t2/p_1_in [7]),
        .I2(\r6/t1/t1/p_0_in [7]),
        .I3(k5b[111]),
        .I4(\r6/t3/t3/p_1_in [7]),
        .I5(\r6/t3/t3/p_0_in [7]),
        .O(\r6/p_0_out [111]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[111]_i_1__5 
       (.I0(\r7/t0/t0/p_0_in [7]),
        .I1(\r7/t2/t2/p_1_in [7]),
        .I2(\r7/t1/t1/p_0_in [7]),
        .I3(k6b[111]),
        .I4(\r7/t3/t3/p_1_in [7]),
        .I5(\r7/t3/t3/p_0_in [7]),
        .O(\r7/p_0_out [111]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[111]_i_1__6 
       (.I0(\r8/t0/t0/p_0_in [7]),
        .I1(\r8/t2/t2/p_1_in [7]),
        .I2(\r8/t1/t1/p_0_in [7]),
        .I3(k7b[111]),
        .I4(\r8/t3/t3/p_1_in [7]),
        .I5(\r8/t3/t3/p_0_in [7]),
        .O(\r8/p_0_out [111]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[111]_i_1__7 
       (.I0(\r9/t0/t0/p_0_in [7]),
        .I1(\r9/t2/t2/p_1_in [7]),
        .I2(\r9/t1/t1/p_0_in [7]),
        .I3(k8b[111]),
        .I4(\r9/t3/t3/p_1_in [7]),
        .I5(\r9/t3/t3/p_0_in [7]),
        .O(\r9/p_0_out [111]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair382" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[111]_i_1__8 
       (.I0(\a10/k0a [15]),
        .I1(\a10/k4a [15]),
        .I2(\rf/p_3_in [15]),
        .O(\rf/p_4_out [111]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[112]_i_1 
       (.I0(\r1/t0/t0/p_0_in [0]),
        .I1(\r1/t2/t2/p_1_in [0]),
        .I2(\r1/t2/t2/p_0_in [0]),
        .I3(\r1/t1/t1/p_1_in [0]),
        .I4(k0b[112]),
        .I5(\r1/t3/t3/p_0_in [0]),
        .O(\r1/p_0_out [112]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[112]_i_1__0 
       (.I0(\r2/t0/t0/p_0_in [0]),
        .I1(\r2/t2/t2/p_1_in [0]),
        .I2(\r2/t2/t2/p_0_in [0]),
        .I3(\r2/t1/t1/p_1_in [0]),
        .I4(k1b[112]),
        .I5(\r2/t3/t3/p_0_in [0]),
        .O(\r2/p_0_out [112]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[112]_i_1__1 
       (.I0(\r3/t0/t0/p_0_in [0]),
        .I1(\r3/t2/t2/p_1_in [0]),
        .I2(\r3/t2/t2/p_0_in [0]),
        .I3(\r3/t1/t1/p_1_in [0]),
        .I4(k2b[112]),
        .I5(\r3/t3/t3/p_0_in [0]),
        .O(\r3/p_0_out [112]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[112]_i_1__2 
       (.I0(\r4/t0/t0/p_0_in [0]),
        .I1(\r4/t2/t2/p_1_in [0]),
        .I2(\r4/t2/t2/p_0_in [0]),
        .I3(\r4/t1/t1/p_1_in [0]),
        .I4(k3b[112]),
        .I5(\r4/t3/t3/p_0_in [0]),
        .O(\r4/p_0_out [112]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[112]_i_1__3 
       (.I0(\r5/t0/t0/p_0_in [0]),
        .I1(\r5/t2/t2/p_1_in [0]),
        .I2(\r5/t2/t2/p_0_in [0]),
        .I3(\r5/t1/t1/p_1_in [0]),
        .I4(k4b[112]),
        .I5(\r5/t3/t3/p_0_in [0]),
        .O(\r5/p_0_out [112]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[112]_i_1__4 
       (.I0(\r6/t0/t0/p_0_in [0]),
        .I1(\r6/t2/t2/p_1_in [0]),
        .I2(\r6/t2/t2/p_0_in [0]),
        .I3(\r6/t1/t1/p_1_in [0]),
        .I4(k5b[112]),
        .I5(\r6/t3/t3/p_0_in [0]),
        .O(\r6/p_0_out [112]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[112]_i_1__5 
       (.I0(\r7/t0/t0/p_0_in [0]),
        .I1(\r7/t2/t2/p_1_in [0]),
        .I2(\r7/t2/t2/p_0_in [0]),
        .I3(\r7/t1/t1/p_1_in [0]),
        .I4(k6b[112]),
        .I5(\r7/t3/t3/p_0_in [0]),
        .O(\r7/p_0_out [112]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[112]_i_1__6 
       (.I0(\r8/t0/t0/p_0_in [0]),
        .I1(\r8/t2/t2/p_1_in [0]),
        .I2(\r8/t2/t2/p_0_in [0]),
        .I3(\r8/t1/t1/p_1_in [0]),
        .I4(k7b[112]),
        .I5(\r8/t3/t3/p_0_in [0]),
        .O(\r8/p_0_out [112]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[112]_i_1__7 
       (.I0(\r9/t0/t0/p_0_in [0]),
        .I1(\r9/t2/t2/p_1_in [0]),
        .I2(\r9/t2/t2/p_0_in [0]),
        .I3(\r9/t1/t1/p_1_in [0]),
        .I4(k8b[112]),
        .I5(\r9/t3/t3/p_0_in [0]),
        .O(\r9/p_0_out [112]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair381" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[112]_i_1__8 
       (.I0(\a10/k0a [16]),
        .I1(\a10/k4a [16]),
        .I2(\rf/p_3_in [16]),
        .O(\rf/p_4_out [112]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[113]_i_1 
       (.I0(\r1/t0/t0/p_0_in [1]),
        .I1(\r1/t2/t2/p_1_in [1]),
        .I2(\r1/t2/t2/p_0_in [1]),
        .I3(\r1/t1/t1/p_1_in [1]),
        .I4(k0b[113]),
        .I5(\r1/t3/t3/p_0_in [1]),
        .O(\r1/p_0_out [113]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[113]_i_1__0 
       (.I0(\r2/t0/t0/p_0_in [1]),
        .I1(\r2/t2/t2/p_1_in [1]),
        .I2(\r2/t2/t2/p_0_in [1]),
        .I3(\r2/t1/t1/p_1_in [1]),
        .I4(k1b[113]),
        .I5(\r2/t3/t3/p_0_in [1]),
        .O(\r2/p_0_out [113]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[113]_i_1__1 
       (.I0(\r3/t0/t0/p_0_in [1]),
        .I1(\r3/t2/t2/p_1_in [1]),
        .I2(\r3/t2/t2/p_0_in [1]),
        .I3(\r3/t1/t1/p_1_in [1]),
        .I4(k2b[113]),
        .I5(\r3/t3/t3/p_0_in [1]),
        .O(\r3/p_0_out [113]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[113]_i_1__2 
       (.I0(\r4/t0/t0/p_0_in [1]),
        .I1(\r4/t2/t2/p_1_in [1]),
        .I2(\r4/t2/t2/p_0_in [1]),
        .I3(\r4/t1/t1/p_1_in [1]),
        .I4(k3b[113]),
        .I5(\r4/t3/t3/p_0_in [1]),
        .O(\r4/p_0_out [113]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[113]_i_1__3 
       (.I0(\r5/t0/t0/p_0_in [1]),
        .I1(\r5/t2/t2/p_1_in [1]),
        .I2(\r5/t2/t2/p_0_in [1]),
        .I3(\r5/t1/t1/p_1_in [1]),
        .I4(k4b[113]),
        .I5(\r5/t3/t3/p_0_in [1]),
        .O(\r5/p_0_out [113]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[113]_i_1__4 
       (.I0(\r6/t0/t0/p_0_in [1]),
        .I1(\r6/t2/t2/p_1_in [1]),
        .I2(\r6/t2/t2/p_0_in [1]),
        .I3(\r6/t1/t1/p_1_in [1]),
        .I4(k5b[113]),
        .I5(\r6/t3/t3/p_0_in [1]),
        .O(\r6/p_0_out [113]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[113]_i_1__5 
       (.I0(\r7/t0/t0/p_0_in [1]),
        .I1(\r7/t2/t2/p_1_in [1]),
        .I2(\r7/t2/t2/p_0_in [1]),
        .I3(\r7/t1/t1/p_1_in [1]),
        .I4(k6b[113]),
        .I5(\r7/t3/t3/p_0_in [1]),
        .O(\r7/p_0_out [113]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[113]_i_1__6 
       (.I0(\r8/t0/t0/p_0_in [1]),
        .I1(\r8/t2/t2/p_1_in [1]),
        .I2(\r8/t2/t2/p_0_in [1]),
        .I3(\r8/t1/t1/p_1_in [1]),
        .I4(k7b[113]),
        .I5(\r8/t3/t3/p_0_in [1]),
        .O(\r8/p_0_out [113]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[113]_i_1__7 
       (.I0(\r9/t0/t0/p_0_in [1]),
        .I1(\r9/t2/t2/p_1_in [1]),
        .I2(\r9/t2/t2/p_0_in [1]),
        .I3(\r9/t1/t1/p_1_in [1]),
        .I4(k8b[113]),
        .I5(\r9/t3/t3/p_0_in [1]),
        .O(\r9/p_0_out [113]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair380" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[113]_i_1__8 
       (.I0(\a10/k0a [17]),
        .I1(\a10/k4a [17]),
        .I2(\rf/p_3_in [17]),
        .O(\rf/p_4_out [113]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[114]_i_1 
       (.I0(\r1/t0/t0/p_0_in [2]),
        .I1(\r1/t2/t2/p_1_in [2]),
        .I2(\r1/t2/t2/p_0_in [2]),
        .I3(\r1/t1/t1/p_1_in [2]),
        .I4(k0b[114]),
        .I5(\r1/t3/t3/p_0_in [2]),
        .O(\r1/p_0_out [114]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[114]_i_1__0 
       (.I0(\r2/t0/t0/p_0_in [2]),
        .I1(\r2/t2/t2/p_1_in [2]),
        .I2(\r2/t2/t2/p_0_in [2]),
        .I3(\r2/t1/t1/p_1_in [2]),
        .I4(k1b[114]),
        .I5(\r2/t3/t3/p_0_in [2]),
        .O(\r2/p_0_out [114]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[114]_i_1__1 
       (.I0(\r3/t0/t0/p_0_in [2]),
        .I1(\r3/t2/t2/p_1_in [2]),
        .I2(\r3/t2/t2/p_0_in [2]),
        .I3(\r3/t1/t1/p_1_in [2]),
        .I4(k2b[114]),
        .I5(\r3/t3/t3/p_0_in [2]),
        .O(\r3/p_0_out [114]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[114]_i_1__2 
       (.I0(\r4/t0/t0/p_0_in [2]),
        .I1(\r4/t2/t2/p_1_in [2]),
        .I2(\r4/t2/t2/p_0_in [2]),
        .I3(\r4/t1/t1/p_1_in [2]),
        .I4(k3b[114]),
        .I5(\r4/t3/t3/p_0_in [2]),
        .O(\r4/p_0_out [114]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[114]_i_1__3 
       (.I0(\r5/t0/t0/p_0_in [2]),
        .I1(\r5/t2/t2/p_1_in [2]),
        .I2(\r5/t2/t2/p_0_in [2]),
        .I3(\r5/t1/t1/p_1_in [2]),
        .I4(k4b[114]),
        .I5(\r5/t3/t3/p_0_in [2]),
        .O(\r5/p_0_out [114]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[114]_i_1__4 
       (.I0(\r6/t0/t0/p_0_in [2]),
        .I1(\r6/t2/t2/p_1_in [2]),
        .I2(\r6/t2/t2/p_0_in [2]),
        .I3(\r6/t1/t1/p_1_in [2]),
        .I4(k5b[114]),
        .I5(\r6/t3/t3/p_0_in [2]),
        .O(\r6/p_0_out [114]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[114]_i_1__5 
       (.I0(\r7/t0/t0/p_0_in [2]),
        .I1(\r7/t2/t2/p_1_in [2]),
        .I2(\r7/t2/t2/p_0_in [2]),
        .I3(\r7/t1/t1/p_1_in [2]),
        .I4(k6b[114]),
        .I5(\r7/t3/t3/p_0_in [2]),
        .O(\r7/p_0_out [114]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[114]_i_1__6 
       (.I0(\r8/t0/t0/p_0_in [2]),
        .I1(\r8/t2/t2/p_1_in [2]),
        .I2(\r8/t2/t2/p_0_in [2]),
        .I3(\r8/t1/t1/p_1_in [2]),
        .I4(k7b[114]),
        .I5(\r8/t3/t3/p_0_in [2]),
        .O(\r8/p_0_out [114]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[114]_i_1__7 
       (.I0(\r9/t0/t0/p_0_in [2]),
        .I1(\r9/t2/t2/p_1_in [2]),
        .I2(\r9/t2/t2/p_0_in [2]),
        .I3(\r9/t1/t1/p_1_in [2]),
        .I4(k8b[114]),
        .I5(\r9/t3/t3/p_0_in [2]),
        .O(\r9/p_0_out [114]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair379" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[114]_i_1__8 
       (.I0(\a10/k0a [18]),
        .I1(\a10/k4a [18]),
        .I2(\rf/p_3_in [18]),
        .O(\rf/p_4_out [114]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[115]_i_1 
       (.I0(\r1/t0/t0/p_0_in [3]),
        .I1(\r1/t2/t2/p_1_in [3]),
        .I2(\r1/t2/t2/p_0_in [3]),
        .I3(\r1/t1/t1/p_1_in [3]),
        .I4(k0b[115]),
        .I5(\r1/t3/t3/p_0_in [3]),
        .O(\r1/p_0_out [115]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[115]_i_1__0 
       (.I0(\r2/t0/t0/p_0_in [3]),
        .I1(\r2/t2/t2/p_1_in [3]),
        .I2(\r2/t2/t2/p_0_in [3]),
        .I3(\r2/t1/t1/p_1_in [3]),
        .I4(k1b[115]),
        .I5(\r2/t3/t3/p_0_in [3]),
        .O(\r2/p_0_out [115]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[115]_i_1__1 
       (.I0(\r3/t0/t0/p_0_in [3]),
        .I1(\r3/t2/t2/p_1_in [3]),
        .I2(\r3/t2/t2/p_0_in [3]),
        .I3(\r3/t1/t1/p_1_in [3]),
        .I4(k2b[115]),
        .I5(\r3/t3/t3/p_0_in [3]),
        .O(\r3/p_0_out [115]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[115]_i_1__2 
       (.I0(\r4/t0/t0/p_0_in [3]),
        .I1(\r4/t2/t2/p_1_in [3]),
        .I2(\r4/t2/t2/p_0_in [3]),
        .I3(\r4/t1/t1/p_1_in [3]),
        .I4(k3b[115]),
        .I5(\r4/t3/t3/p_0_in [3]),
        .O(\r4/p_0_out [115]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[115]_i_1__3 
       (.I0(\r5/t0/t0/p_0_in [3]),
        .I1(\r5/t2/t2/p_1_in [3]),
        .I2(\r5/t2/t2/p_0_in [3]),
        .I3(\r5/t1/t1/p_1_in [3]),
        .I4(k4b[115]),
        .I5(\r5/t3/t3/p_0_in [3]),
        .O(\r5/p_0_out [115]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[115]_i_1__4 
       (.I0(\r6/t0/t0/p_0_in [3]),
        .I1(\r6/t2/t2/p_1_in [3]),
        .I2(\r6/t2/t2/p_0_in [3]),
        .I3(\r6/t1/t1/p_1_in [3]),
        .I4(k5b[115]),
        .I5(\r6/t3/t3/p_0_in [3]),
        .O(\r6/p_0_out [115]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[115]_i_1__5 
       (.I0(\r7/t0/t0/p_0_in [3]),
        .I1(\r7/t2/t2/p_1_in [3]),
        .I2(\r7/t2/t2/p_0_in [3]),
        .I3(\r7/t1/t1/p_1_in [3]),
        .I4(k6b[115]),
        .I5(\r7/t3/t3/p_0_in [3]),
        .O(\r7/p_0_out [115]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[115]_i_1__6 
       (.I0(\r8/t0/t0/p_0_in [3]),
        .I1(\r8/t2/t2/p_1_in [3]),
        .I2(\r8/t2/t2/p_0_in [3]),
        .I3(\r8/t1/t1/p_1_in [3]),
        .I4(k7b[115]),
        .I5(\r8/t3/t3/p_0_in [3]),
        .O(\r8/p_0_out [115]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[115]_i_1__7 
       (.I0(\r9/t0/t0/p_0_in [3]),
        .I1(\r9/t2/t2/p_1_in [3]),
        .I2(\r9/t2/t2/p_0_in [3]),
        .I3(\r9/t1/t1/p_1_in [3]),
        .I4(k8b[115]),
        .I5(\r9/t3/t3/p_0_in [3]),
        .O(\r9/p_0_out [115]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair378" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[115]_i_1__8 
       (.I0(\a10/k0a [19]),
        .I1(\a10/k4a [19]),
        .I2(\rf/p_3_in [19]),
        .O(\rf/p_4_out [115]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[116]_i_1 
       (.I0(\r1/t0/t0/p_0_in [4]),
        .I1(\r1/t2/t2/p_1_in [4]),
        .I2(\r1/t2/t2/p_0_in [4]),
        .I3(\r1/t1/t1/p_1_in [4]),
        .I4(k0b[116]),
        .I5(\r1/t3/t3/p_0_in [4]),
        .O(\r1/p_0_out [116]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[116]_i_1__0 
       (.I0(\r2/t0/t0/p_0_in [4]),
        .I1(\r2/t2/t2/p_1_in [4]),
        .I2(\r2/t2/t2/p_0_in [4]),
        .I3(\r2/t1/t1/p_1_in [4]),
        .I4(k1b[116]),
        .I5(\r2/t3/t3/p_0_in [4]),
        .O(\r2/p_0_out [116]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[116]_i_1__1 
       (.I0(\r3/t0/t0/p_0_in [4]),
        .I1(\r3/t2/t2/p_1_in [4]),
        .I2(\r3/t2/t2/p_0_in [4]),
        .I3(\r3/t1/t1/p_1_in [4]),
        .I4(k2b[116]),
        .I5(\r3/t3/t3/p_0_in [4]),
        .O(\r3/p_0_out [116]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[116]_i_1__2 
       (.I0(\r4/t0/t0/p_0_in [4]),
        .I1(\r4/t2/t2/p_1_in [4]),
        .I2(\r4/t2/t2/p_0_in [4]),
        .I3(\r4/t1/t1/p_1_in [4]),
        .I4(k3b[116]),
        .I5(\r4/t3/t3/p_0_in [4]),
        .O(\r4/p_0_out [116]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[116]_i_1__3 
       (.I0(\r5/t0/t0/p_0_in [4]),
        .I1(\r5/t2/t2/p_1_in [4]),
        .I2(\r5/t2/t2/p_0_in [4]),
        .I3(\r5/t1/t1/p_1_in [4]),
        .I4(k4b[116]),
        .I5(\r5/t3/t3/p_0_in [4]),
        .O(\r5/p_0_out [116]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[116]_i_1__4 
       (.I0(\r6/t0/t0/p_0_in [4]),
        .I1(\r6/t2/t2/p_1_in [4]),
        .I2(\r6/t2/t2/p_0_in [4]),
        .I3(\r6/t1/t1/p_1_in [4]),
        .I4(k5b[116]),
        .I5(\r6/t3/t3/p_0_in [4]),
        .O(\r6/p_0_out [116]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[116]_i_1__5 
       (.I0(\r7/t0/t0/p_0_in [4]),
        .I1(\r7/t2/t2/p_1_in [4]),
        .I2(\r7/t2/t2/p_0_in [4]),
        .I3(\r7/t1/t1/p_1_in [4]),
        .I4(k6b[116]),
        .I5(\r7/t3/t3/p_0_in [4]),
        .O(\r7/p_0_out [116]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[116]_i_1__6 
       (.I0(\r8/t0/t0/p_0_in [4]),
        .I1(\r8/t2/t2/p_1_in [4]),
        .I2(\r8/t2/t2/p_0_in [4]),
        .I3(\r8/t1/t1/p_1_in [4]),
        .I4(k7b[116]),
        .I5(\r8/t3/t3/p_0_in [4]),
        .O(\r8/p_0_out [116]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[116]_i_1__7 
       (.I0(\r9/t0/t0/p_0_in [4]),
        .I1(\r9/t2/t2/p_1_in [4]),
        .I2(\r9/t2/t2/p_0_in [4]),
        .I3(\r9/t1/t1/p_1_in [4]),
        .I4(k8b[116]),
        .I5(\r9/t3/t3/p_0_in [4]),
        .O(\r9/p_0_out [116]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair377" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[116]_i_1__8 
       (.I0(\a10/k0a [20]),
        .I1(\a10/k4a [20]),
        .I2(\rf/p_3_in [20]),
        .O(\rf/p_4_out [116]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[117]_i_1 
       (.I0(\r1/t0/t0/p_0_in [5]),
        .I1(\r1/t2/t2/p_1_in [5]),
        .I2(\r1/t2/t2/p_0_in [5]),
        .I3(\r1/t1/t1/p_1_in [5]),
        .I4(k0b[117]),
        .I5(\r1/t3/t3/p_0_in [5]),
        .O(\r1/p_0_out [117]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[117]_i_1__0 
       (.I0(\r2/t0/t0/p_0_in [5]),
        .I1(\r2/t2/t2/p_1_in [5]),
        .I2(\r2/t2/t2/p_0_in [5]),
        .I3(\r2/t1/t1/p_1_in [5]),
        .I4(k1b[117]),
        .I5(\r2/t3/t3/p_0_in [5]),
        .O(\r2/p_0_out [117]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[117]_i_1__1 
       (.I0(\r3/t0/t0/p_0_in [5]),
        .I1(\r3/t2/t2/p_1_in [5]),
        .I2(\r3/t2/t2/p_0_in [5]),
        .I3(\r3/t1/t1/p_1_in [5]),
        .I4(k2b[117]),
        .I5(\r3/t3/t3/p_0_in [5]),
        .O(\r3/p_0_out [117]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[117]_i_1__2 
       (.I0(\r4/t0/t0/p_0_in [5]),
        .I1(\r4/t2/t2/p_1_in [5]),
        .I2(\r4/t2/t2/p_0_in [5]),
        .I3(\r4/t1/t1/p_1_in [5]),
        .I4(k3b[117]),
        .I5(\r4/t3/t3/p_0_in [5]),
        .O(\r4/p_0_out [117]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[117]_i_1__3 
       (.I0(\r5/t0/t0/p_0_in [5]),
        .I1(\r5/t2/t2/p_1_in [5]),
        .I2(\r5/t2/t2/p_0_in [5]),
        .I3(\r5/t1/t1/p_1_in [5]),
        .I4(k4b[117]),
        .I5(\r5/t3/t3/p_0_in [5]),
        .O(\r5/p_0_out [117]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[117]_i_1__4 
       (.I0(\r6/t0/t0/p_0_in [5]),
        .I1(\r6/t2/t2/p_1_in [5]),
        .I2(\r6/t2/t2/p_0_in [5]),
        .I3(\r6/t1/t1/p_1_in [5]),
        .I4(k5b[117]),
        .I5(\r6/t3/t3/p_0_in [5]),
        .O(\r6/p_0_out [117]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[117]_i_1__5 
       (.I0(\r7/t0/t0/p_0_in [5]),
        .I1(\r7/t2/t2/p_1_in [5]),
        .I2(\r7/t2/t2/p_0_in [5]),
        .I3(\r7/t1/t1/p_1_in [5]),
        .I4(k6b[117]),
        .I5(\r7/t3/t3/p_0_in [5]),
        .O(\r7/p_0_out [117]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[117]_i_1__6 
       (.I0(\r8/t0/t0/p_0_in [5]),
        .I1(\r8/t2/t2/p_1_in [5]),
        .I2(\r8/t2/t2/p_0_in [5]),
        .I3(\r8/t1/t1/p_1_in [5]),
        .I4(k7b[117]),
        .I5(\r8/t3/t3/p_0_in [5]),
        .O(\r8/p_0_out [117]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[117]_i_1__7 
       (.I0(\r9/t0/t0/p_0_in [5]),
        .I1(\r9/t2/t2/p_1_in [5]),
        .I2(\r9/t2/t2/p_0_in [5]),
        .I3(\r9/t1/t1/p_1_in [5]),
        .I4(k8b[117]),
        .I5(\r9/t3/t3/p_0_in [5]),
        .O(\r9/p_0_out [117]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair376" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[117]_i_1__8 
       (.I0(\a10/k0a [21]),
        .I1(\a10/k4a [21]),
        .I2(\rf/p_3_in [21]),
        .O(\rf/p_4_out [117]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[118]_i_1 
       (.I0(\r1/t0/t0/p_0_in [6]),
        .I1(\r1/t2/t2/p_1_in [6]),
        .I2(\r1/t2/t2/p_0_in [6]),
        .I3(\r1/t1/t1/p_1_in [6]),
        .I4(k0b[118]),
        .I5(\r1/t3/t3/p_0_in [6]),
        .O(\r1/p_0_out [118]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[118]_i_1__0 
       (.I0(\r2/t0/t0/p_0_in [6]),
        .I1(\r2/t2/t2/p_1_in [6]),
        .I2(\r2/t2/t2/p_0_in [6]),
        .I3(\r2/t1/t1/p_1_in [6]),
        .I4(k1b[118]),
        .I5(\r2/t3/t3/p_0_in [6]),
        .O(\r2/p_0_out [118]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[118]_i_1__1 
       (.I0(\r3/t0/t0/p_0_in [6]),
        .I1(\r3/t2/t2/p_1_in [6]),
        .I2(\r3/t2/t2/p_0_in [6]),
        .I3(\r3/t1/t1/p_1_in [6]),
        .I4(k2b[118]),
        .I5(\r3/t3/t3/p_0_in [6]),
        .O(\r3/p_0_out [118]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[118]_i_1__2 
       (.I0(\r4/t0/t0/p_0_in [6]),
        .I1(\r4/t2/t2/p_1_in [6]),
        .I2(\r4/t2/t2/p_0_in [6]),
        .I3(\r4/t1/t1/p_1_in [6]),
        .I4(k3b[118]),
        .I5(\r4/t3/t3/p_0_in [6]),
        .O(\r4/p_0_out [118]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[118]_i_1__3 
       (.I0(\r5/t0/t0/p_0_in [6]),
        .I1(\r5/t2/t2/p_1_in [6]),
        .I2(\r5/t2/t2/p_0_in [6]),
        .I3(\r5/t1/t1/p_1_in [6]),
        .I4(k4b[118]),
        .I5(\r5/t3/t3/p_0_in [6]),
        .O(\r5/p_0_out [118]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[118]_i_1__4 
       (.I0(\r6/t0/t0/p_0_in [6]),
        .I1(\r6/t2/t2/p_1_in [6]),
        .I2(\r6/t2/t2/p_0_in [6]),
        .I3(\r6/t1/t1/p_1_in [6]),
        .I4(k5b[118]),
        .I5(\r6/t3/t3/p_0_in [6]),
        .O(\r6/p_0_out [118]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[118]_i_1__5 
       (.I0(\r7/t0/t0/p_0_in [6]),
        .I1(\r7/t2/t2/p_1_in [6]),
        .I2(\r7/t2/t2/p_0_in [6]),
        .I3(\r7/t1/t1/p_1_in [6]),
        .I4(k6b[118]),
        .I5(\r7/t3/t3/p_0_in [6]),
        .O(\r7/p_0_out [118]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[118]_i_1__6 
       (.I0(\r8/t0/t0/p_0_in [6]),
        .I1(\r8/t2/t2/p_1_in [6]),
        .I2(\r8/t2/t2/p_0_in [6]),
        .I3(\r8/t1/t1/p_1_in [6]),
        .I4(k7b[118]),
        .I5(\r8/t3/t3/p_0_in [6]),
        .O(\r8/p_0_out [118]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[118]_i_1__7 
       (.I0(\r9/t0/t0/p_0_in [6]),
        .I1(\r9/t2/t2/p_1_in [6]),
        .I2(\r9/t2/t2/p_0_in [6]),
        .I3(\r9/t1/t1/p_1_in [6]),
        .I4(k8b[118]),
        .I5(\r9/t3/t3/p_0_in [6]),
        .O(\r9/p_0_out [118]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair375" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[118]_i_1__8 
       (.I0(\a10/k0a [22]),
        .I1(\a10/k4a [22]),
        .I2(\rf/p_3_in [22]),
        .O(\rf/p_4_out [118]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[119]_i_1 
       (.I0(\r1/t0/t0/p_0_in [7]),
        .I1(\r1/t2/t2/p_1_in [7]),
        .I2(\r1/t2/t2/p_0_in [7]),
        .I3(\r1/t1/t1/p_1_in [7]),
        .I4(k0b[119]),
        .I5(\r1/t3/t3/p_0_in [7]),
        .O(\r1/p_0_out [119]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[119]_i_1__0 
       (.I0(\r2/t0/t0/p_0_in [7]),
        .I1(\r2/t2/t2/p_1_in [7]),
        .I2(\r2/t2/t2/p_0_in [7]),
        .I3(\r2/t1/t1/p_1_in [7]),
        .I4(k1b[119]),
        .I5(\r2/t3/t3/p_0_in [7]),
        .O(\r2/p_0_out [119]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[119]_i_1__1 
       (.I0(\r3/t0/t0/p_0_in [7]),
        .I1(\r3/t2/t2/p_1_in [7]),
        .I2(\r3/t2/t2/p_0_in [7]),
        .I3(\r3/t1/t1/p_1_in [7]),
        .I4(k2b[119]),
        .I5(\r3/t3/t3/p_0_in [7]),
        .O(\r3/p_0_out [119]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[119]_i_1__2 
       (.I0(\r4/t0/t0/p_0_in [7]),
        .I1(\r4/t2/t2/p_1_in [7]),
        .I2(\r4/t2/t2/p_0_in [7]),
        .I3(\r4/t1/t1/p_1_in [7]),
        .I4(k3b[119]),
        .I5(\r4/t3/t3/p_0_in [7]),
        .O(\r4/p_0_out [119]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[119]_i_1__3 
       (.I0(\r5/t0/t0/p_0_in [7]),
        .I1(\r5/t2/t2/p_1_in [7]),
        .I2(\r5/t2/t2/p_0_in [7]),
        .I3(\r5/t1/t1/p_1_in [7]),
        .I4(k4b[119]),
        .I5(\r5/t3/t3/p_0_in [7]),
        .O(\r5/p_0_out [119]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[119]_i_1__4 
       (.I0(\r6/t0/t0/p_0_in [7]),
        .I1(\r6/t2/t2/p_1_in [7]),
        .I2(\r6/t2/t2/p_0_in [7]),
        .I3(\r6/t1/t1/p_1_in [7]),
        .I4(k5b[119]),
        .I5(\r6/t3/t3/p_0_in [7]),
        .O(\r6/p_0_out [119]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[119]_i_1__5 
       (.I0(\r7/t0/t0/p_0_in [7]),
        .I1(\r7/t2/t2/p_1_in [7]),
        .I2(\r7/t2/t2/p_0_in [7]),
        .I3(\r7/t1/t1/p_1_in [7]),
        .I4(k6b[119]),
        .I5(\r7/t3/t3/p_0_in [7]),
        .O(\r7/p_0_out [119]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[119]_i_1__6 
       (.I0(\r8/t0/t0/p_0_in [7]),
        .I1(\r8/t2/t2/p_1_in [7]),
        .I2(\r8/t2/t2/p_0_in [7]),
        .I3(\r8/t1/t1/p_1_in [7]),
        .I4(k7b[119]),
        .I5(\r8/t3/t3/p_0_in [7]),
        .O(\r8/p_0_out [119]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[119]_i_1__7 
       (.I0(\r9/t0/t0/p_0_in [7]),
        .I1(\r9/t2/t2/p_1_in [7]),
        .I2(\r9/t2/t2/p_0_in [7]),
        .I3(\r9/t1/t1/p_1_in [7]),
        .I4(k8b[119]),
        .I5(\r9/t3/t3/p_0_in [7]),
        .O(\r9/p_0_out [119]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair360" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[119]_i_1__8 
       (.I0(\a10/k0a [23]),
        .I1(\a10/k4a [23]),
        .I2(\rf/p_3_in [23]),
        .O(\rf/p_4_out [119]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[11]_i_1 
       (.I0(\r1/t0/t1/p_0_in [3]),
        .I1(\r1/t2/t3/p_1_in [3]),
        .I2(\r1/t2/t3/p_0_in [3]),
        .I3(\r1/t1/t2/p_1_in [3]),
        .I4(k0b[11]),
        .I5(\r1/t3/t0/p_0_in [3]),
        .O(\r1/p_0_out [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[11]_i_1__0 
       (.I0(\r2/t0/t1/p_0_in [3]),
        .I1(\r2/t2/t3/p_1_in [3]),
        .I2(\r2/t2/t3/p_0_in [3]),
        .I3(\r2/t1/t2/p_1_in [3]),
        .I4(k1b[11]),
        .I5(\r2/t3/t0/p_0_in [3]),
        .O(\r2/p_0_out [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[11]_i_1__1 
       (.I0(\r3/t0/t1/p_0_in [3]),
        .I1(\r3/t2/t3/p_1_in [3]),
        .I2(\r3/t2/t3/p_0_in [3]),
        .I3(\r3/t1/t2/p_1_in [3]),
        .I4(k2b[11]),
        .I5(\r3/t3/t0/p_0_in [3]),
        .O(\r3/p_0_out [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[11]_i_1__2 
       (.I0(\r4/t0/t1/p_0_in [3]),
        .I1(\r4/t2/t3/p_1_in [3]),
        .I2(\r4/t2/t3/p_0_in [3]),
        .I3(\r4/t1/t2/p_1_in [3]),
        .I4(k3b[11]),
        .I5(\r4/t3/t0/p_0_in [3]),
        .O(\r4/p_0_out [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[11]_i_1__3 
       (.I0(\r5/t0/t1/p_0_in [3]),
        .I1(\r5/t2/t3/p_1_in [3]),
        .I2(\r5/t2/t3/p_0_in [3]),
        .I3(\r5/t1/t2/p_1_in [3]),
        .I4(k4b[11]),
        .I5(\r5/t3/t0/p_0_in [3]),
        .O(\r5/p_0_out [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[11]_i_1__4 
       (.I0(\r6/t0/t1/p_0_in [3]),
        .I1(\r6/t2/t3/p_1_in [3]),
        .I2(\r6/t2/t3/p_0_in [3]),
        .I3(\r6/t1/t2/p_1_in [3]),
        .I4(k5b[11]),
        .I5(\r6/t3/t0/p_0_in [3]),
        .O(\r6/p_0_out [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[11]_i_1__5 
       (.I0(\r7/t0/t1/p_0_in [3]),
        .I1(\r7/t2/t3/p_1_in [3]),
        .I2(\r7/t2/t3/p_0_in [3]),
        .I3(\r7/t1/t2/p_1_in [3]),
        .I4(k6b[11]),
        .I5(\r7/t3/t0/p_0_in [3]),
        .O(\r7/p_0_out [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[11]_i_1__6 
       (.I0(\r8/t0/t1/p_0_in [3]),
        .I1(\r8/t2/t3/p_1_in [3]),
        .I2(\r8/t2/t3/p_0_in [3]),
        .I3(\r8/t1/t2/p_1_in [3]),
        .I4(k7b[11]),
        .I5(\r8/t3/t0/p_0_in [3]),
        .O(\r8/p_0_out [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[11]_i_1__7 
       (.I0(\r9/t0/t1/p_0_in [3]),
        .I1(\r9/t2/t3/p_1_in [3]),
        .I2(\r9/t2/t3/p_0_in [3]),
        .I3(\r9/t1/t2/p_1_in [3]),
        .I4(k8b[11]),
        .I5(\r9/t3/t0/p_0_in [3]),
        .O(\r9/p_0_out [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair331" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[11]_i_1__8 
       (.I0(\a10/k3a [11]),
        .I1(\a10/k4a [11]),
        .I2(\rf/p_0_in [11]),
        .O(\rf/p_4_out [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[120]_i_1 
       (.I0(\r1/t0/t0/p_1_in [0]),
        .I1(\r1/t2/t2/p_0_in [0]),
        .I2(\r1/t1/t1/p_1_in [0]),
        .I3(\r1/t1/t1/p_0_in [0]),
        .I4(k0b[120]),
        .I5(\r1/t3/t3/p_0_in [0]),
        .O(\r1/p_0_out [120]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[120]_i_1__0 
       (.I0(\r2/t0/t0/p_1_in [0]),
        .I1(\r2/t2/t2/p_0_in [0]),
        .I2(\r2/t1/t1/p_1_in [0]),
        .I3(\r2/t1/t1/p_0_in [0]),
        .I4(k1b[120]),
        .I5(\r2/t3/t3/p_0_in [0]),
        .O(\r2/p_0_out [120]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[120]_i_1__1 
       (.I0(\r3/t0/t0/p_1_in [0]),
        .I1(\r3/t2/t2/p_0_in [0]),
        .I2(\r3/t1/t1/p_1_in [0]),
        .I3(\r3/t1/t1/p_0_in [0]),
        .I4(k2b[120]),
        .I5(\r3/t3/t3/p_0_in [0]),
        .O(\r3/p_0_out [120]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[120]_i_1__2 
       (.I0(\r4/t0/t0/p_1_in [0]),
        .I1(\r4/t2/t2/p_0_in [0]),
        .I2(\r4/t1/t1/p_1_in [0]),
        .I3(\r4/t1/t1/p_0_in [0]),
        .I4(k3b[120]),
        .I5(\r4/t3/t3/p_0_in [0]),
        .O(\r4/p_0_out [120]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[120]_i_1__3 
       (.I0(\r5/t0/t0/p_1_in [0]),
        .I1(\r5/t2/t2/p_0_in [0]),
        .I2(\r5/t1/t1/p_1_in [0]),
        .I3(\r5/t1/t1/p_0_in [0]),
        .I4(k4b[120]),
        .I5(\r5/t3/t3/p_0_in [0]),
        .O(\r5/p_0_out [120]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[120]_i_1__4 
       (.I0(\r6/t0/t0/p_1_in [0]),
        .I1(\r6/t2/t2/p_0_in [0]),
        .I2(\r6/t1/t1/p_1_in [0]),
        .I3(\r6/t1/t1/p_0_in [0]),
        .I4(k5b[120]),
        .I5(\r6/t3/t3/p_0_in [0]),
        .O(\r6/p_0_out [120]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[120]_i_1__5 
       (.I0(\r7/t0/t0/p_1_in [0]),
        .I1(\r7/t2/t2/p_0_in [0]),
        .I2(\r7/t1/t1/p_1_in [0]),
        .I3(\r7/t1/t1/p_0_in [0]),
        .I4(k6b[120]),
        .I5(\r7/t3/t3/p_0_in [0]),
        .O(\r7/p_0_out [120]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[120]_i_1__6 
       (.I0(\r8/t0/t0/p_1_in [0]),
        .I1(\r8/t2/t2/p_0_in [0]),
        .I2(\r8/t1/t1/p_1_in [0]),
        .I3(\r8/t1/t1/p_0_in [0]),
        .I4(k7b[120]),
        .I5(\r8/t3/t3/p_0_in [0]),
        .O(\r8/p_0_out [120]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[120]_i_1__7 
       (.I0(\r9/t0/t0/p_1_in [0]),
        .I1(\r9/t2/t2/p_0_in [0]),
        .I2(\r9/t1/t1/p_1_in [0]),
        .I3(\r9/t1/t1/p_0_in [0]),
        .I4(k8b[120]),
        .I5(\r9/t3/t3/p_0_in [0]),
        .O(\r9/p_0_out [120]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair325" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[120]_i_1__8 
       (.I0(\a10/k0a [24]),
        .I1(\a10/k4a [24]),
        .I2(\rf/p_3_in [24]),
        .O(\rf/p_4_out [120]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[121]_i_1 
       (.I0(\r1/t0/t0/p_1_in [1]),
        .I1(\r1/t2/t2/p_0_in [1]),
        .I2(\r1/t1/t1/p_1_in [1]),
        .I3(\r1/t1/t1/p_0_in [1]),
        .I4(k0b[121]),
        .I5(\r1/t3/t3/p_0_in [1]),
        .O(\r1/p_0_out [121]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[121]_i_1__0 
       (.I0(\r2/t0/t0/p_1_in [1]),
        .I1(\r2/t2/t2/p_0_in [1]),
        .I2(\r2/t1/t1/p_1_in [1]),
        .I3(\r2/t1/t1/p_0_in [1]),
        .I4(k1b[121]),
        .I5(\r2/t3/t3/p_0_in [1]),
        .O(\r2/p_0_out [121]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[121]_i_1__1 
       (.I0(\r3/t0/t0/p_1_in [1]),
        .I1(\r3/t2/t2/p_0_in [1]),
        .I2(\r3/t1/t1/p_1_in [1]),
        .I3(\r3/t1/t1/p_0_in [1]),
        .I4(k2b[121]),
        .I5(\r3/t3/t3/p_0_in [1]),
        .O(\r3/p_0_out [121]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[121]_i_1__2 
       (.I0(\r4/t0/t0/p_1_in [1]),
        .I1(\r4/t2/t2/p_0_in [1]),
        .I2(\r4/t1/t1/p_1_in [1]),
        .I3(\r4/t1/t1/p_0_in [1]),
        .I4(k3b[121]),
        .I5(\r4/t3/t3/p_0_in [1]),
        .O(\r4/p_0_out [121]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[121]_i_1__3 
       (.I0(\r5/t0/t0/p_1_in [1]),
        .I1(\r5/t2/t2/p_0_in [1]),
        .I2(\r5/t1/t1/p_1_in [1]),
        .I3(\r5/t1/t1/p_0_in [1]),
        .I4(k4b[121]),
        .I5(\r5/t3/t3/p_0_in [1]),
        .O(\r5/p_0_out [121]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[121]_i_1__4 
       (.I0(\r6/t0/t0/p_1_in [1]),
        .I1(\r6/t2/t2/p_0_in [1]),
        .I2(\r6/t1/t1/p_1_in [1]),
        .I3(\r6/t1/t1/p_0_in [1]),
        .I4(k5b[121]),
        .I5(\r6/t3/t3/p_0_in [1]),
        .O(\r6/p_0_out [121]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[121]_i_1__5 
       (.I0(\r7/t0/t0/p_1_in [1]),
        .I1(\r7/t2/t2/p_0_in [1]),
        .I2(\r7/t1/t1/p_1_in [1]),
        .I3(\r7/t1/t1/p_0_in [1]),
        .I4(k6b[121]),
        .I5(\r7/t3/t3/p_0_in [1]),
        .O(\r7/p_0_out [121]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[121]_i_1__6 
       (.I0(\r8/t0/t0/p_1_in [1]),
        .I1(\r8/t2/t2/p_0_in [1]),
        .I2(\r8/t1/t1/p_1_in [1]),
        .I3(\r8/t1/t1/p_0_in [1]),
        .I4(k7b[121]),
        .I5(\r8/t3/t3/p_0_in [1]),
        .O(\r8/p_0_out [121]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[121]_i_1__7 
       (.I0(\r9/t0/t0/p_1_in [1]),
        .I1(\r9/t2/t2/p_0_in [1]),
        .I2(\r9/t1/t1/p_1_in [1]),
        .I3(\r9/t1/t1/p_0_in [1]),
        .I4(k8b[121]),
        .I5(\r9/t3/t3/p_0_in [1]),
        .O(\r9/p_0_out [121]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair322" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[121]_i_1__8 
       (.I0(\a10/k0a [25]),
        .I1(\a10/k4a [25]),
        .I2(\rf/p_3_in [25]),
        .O(\rf/p_4_out [121]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[122]_i_1 
       (.I0(\r1/t0/t0/p_1_in [2]),
        .I1(\r1/t2/t2/p_0_in [2]),
        .I2(\r1/t1/t1/p_1_in [2]),
        .I3(\r1/t1/t1/p_0_in [2]),
        .I4(k0b[122]),
        .I5(\r1/t3/t3/p_0_in [2]),
        .O(\r1/p_0_out [122]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[122]_i_1__0 
       (.I0(\r2/t0/t0/p_1_in [2]),
        .I1(\r2/t2/t2/p_0_in [2]),
        .I2(\r2/t1/t1/p_1_in [2]),
        .I3(\r2/t1/t1/p_0_in [2]),
        .I4(k1b[122]),
        .I5(\r2/t3/t3/p_0_in [2]),
        .O(\r2/p_0_out [122]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[122]_i_1__1 
       (.I0(\r3/t0/t0/p_1_in [2]),
        .I1(\r3/t2/t2/p_0_in [2]),
        .I2(\r3/t1/t1/p_1_in [2]),
        .I3(\r3/t1/t1/p_0_in [2]),
        .I4(k2b[122]),
        .I5(\r3/t3/t3/p_0_in [2]),
        .O(\r3/p_0_out [122]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[122]_i_1__2 
       (.I0(\r4/t0/t0/p_1_in [2]),
        .I1(\r4/t2/t2/p_0_in [2]),
        .I2(\r4/t1/t1/p_1_in [2]),
        .I3(\r4/t1/t1/p_0_in [2]),
        .I4(k3b[122]),
        .I5(\r4/t3/t3/p_0_in [2]),
        .O(\r4/p_0_out [122]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[122]_i_1__3 
       (.I0(\r5/t0/t0/p_1_in [2]),
        .I1(\r5/t2/t2/p_0_in [2]),
        .I2(\r5/t1/t1/p_1_in [2]),
        .I3(\r5/t1/t1/p_0_in [2]),
        .I4(k4b[122]),
        .I5(\r5/t3/t3/p_0_in [2]),
        .O(\r5/p_0_out [122]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[122]_i_1__4 
       (.I0(\r6/t0/t0/p_1_in [2]),
        .I1(\r6/t2/t2/p_0_in [2]),
        .I2(\r6/t1/t1/p_1_in [2]),
        .I3(\r6/t1/t1/p_0_in [2]),
        .I4(k5b[122]),
        .I5(\r6/t3/t3/p_0_in [2]),
        .O(\r6/p_0_out [122]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[122]_i_1__5 
       (.I0(\r7/t0/t0/p_1_in [2]),
        .I1(\r7/t2/t2/p_0_in [2]),
        .I2(\r7/t1/t1/p_1_in [2]),
        .I3(\r7/t1/t1/p_0_in [2]),
        .I4(k6b[122]),
        .I5(\r7/t3/t3/p_0_in [2]),
        .O(\r7/p_0_out [122]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[122]_i_1__6 
       (.I0(\r8/t0/t0/p_1_in [2]),
        .I1(\r8/t2/t2/p_0_in [2]),
        .I2(\r8/t1/t1/p_1_in [2]),
        .I3(\r8/t1/t1/p_0_in [2]),
        .I4(k7b[122]),
        .I5(\r8/t3/t3/p_0_in [2]),
        .O(\r8/p_0_out [122]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[122]_i_1__7 
       (.I0(\r9/t0/t0/p_1_in [2]),
        .I1(\r9/t2/t2/p_0_in [2]),
        .I2(\r9/t1/t1/p_1_in [2]),
        .I3(\r9/t1/t1/p_0_in [2]),
        .I4(k8b[122]),
        .I5(\r9/t3/t3/p_0_in [2]),
        .O(\r9/p_0_out [122]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair327" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[122]_i_1__8 
       (.I0(\a10/k0a [26]),
        .I1(\a10/k4a [26]),
        .I2(\rf/p_3_in [26]),
        .O(\rf/p_4_out [122]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[123]_i_1 
       (.I0(\r1/t0/t0/p_1_in [3]),
        .I1(\r1/t2/t2/p_0_in [3]),
        .I2(\r1/t1/t1/p_1_in [3]),
        .I3(\r1/t1/t1/p_0_in [3]),
        .I4(k0b[123]),
        .I5(\r1/t3/t3/p_0_in [3]),
        .O(\r1/p_0_out [123]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[123]_i_1__0 
       (.I0(\r2/t0/t0/p_1_in [3]),
        .I1(\r2/t2/t2/p_0_in [3]),
        .I2(\r2/t1/t1/p_1_in [3]),
        .I3(\r2/t1/t1/p_0_in [3]),
        .I4(k1b[123]),
        .I5(\r2/t3/t3/p_0_in [3]),
        .O(\r2/p_0_out [123]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[123]_i_1__1 
       (.I0(\r3/t0/t0/p_1_in [3]),
        .I1(\r3/t2/t2/p_0_in [3]),
        .I2(\r3/t1/t1/p_1_in [3]),
        .I3(\r3/t1/t1/p_0_in [3]),
        .I4(k2b[123]),
        .I5(\r3/t3/t3/p_0_in [3]),
        .O(\r3/p_0_out [123]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[123]_i_1__2 
       (.I0(\r4/t0/t0/p_1_in [3]),
        .I1(\r4/t2/t2/p_0_in [3]),
        .I2(\r4/t1/t1/p_1_in [3]),
        .I3(\r4/t1/t1/p_0_in [3]),
        .I4(k3b[123]),
        .I5(\r4/t3/t3/p_0_in [3]),
        .O(\r4/p_0_out [123]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[123]_i_1__3 
       (.I0(\r5/t0/t0/p_1_in [3]),
        .I1(\r5/t2/t2/p_0_in [3]),
        .I2(\r5/t1/t1/p_1_in [3]),
        .I3(\r5/t1/t1/p_0_in [3]),
        .I4(k4b[123]),
        .I5(\r5/t3/t3/p_0_in [3]),
        .O(\r5/p_0_out [123]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[123]_i_1__4 
       (.I0(\r6/t0/t0/p_1_in [3]),
        .I1(\r6/t2/t2/p_0_in [3]),
        .I2(\r6/t1/t1/p_1_in [3]),
        .I3(\r6/t1/t1/p_0_in [3]),
        .I4(k5b[123]),
        .I5(\r6/t3/t3/p_0_in [3]),
        .O(\r6/p_0_out [123]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[123]_i_1__5 
       (.I0(\r7/t0/t0/p_1_in [3]),
        .I1(\r7/t2/t2/p_0_in [3]),
        .I2(\r7/t1/t1/p_1_in [3]),
        .I3(\r7/t1/t1/p_0_in [3]),
        .I4(k6b[123]),
        .I5(\r7/t3/t3/p_0_in [3]),
        .O(\r7/p_0_out [123]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[123]_i_1__6 
       (.I0(\r8/t0/t0/p_1_in [3]),
        .I1(\r8/t2/t2/p_0_in [3]),
        .I2(\r8/t1/t1/p_1_in [3]),
        .I3(\r8/t1/t1/p_0_in [3]),
        .I4(k7b[123]),
        .I5(\r8/t3/t3/p_0_in [3]),
        .O(\r8/p_0_out [123]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[123]_i_1__7 
       (.I0(\r9/t0/t0/p_1_in [3]),
        .I1(\r9/t2/t2/p_0_in [3]),
        .I2(\r9/t1/t1/p_1_in [3]),
        .I3(\r9/t1/t1/p_0_in [3]),
        .I4(k8b[123]),
        .I5(\r9/t3/t3/p_0_in [3]),
        .O(\r9/p_0_out [123]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair326" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[123]_i_1__8 
       (.I0(\a10/k0a [27]),
        .I1(\a10/k4a [27]),
        .I2(\rf/p_3_in [27]),
        .O(\rf/p_4_out [123]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[124]_i_1 
       (.I0(\r1/t0/t0/p_1_in [4]),
        .I1(\r1/t2/t2/p_0_in [4]),
        .I2(\r1/t1/t1/p_1_in [4]),
        .I3(\r1/t1/t1/p_0_in [4]),
        .I4(k0b[124]),
        .I5(\r1/t3/t3/p_0_in [4]),
        .O(\r1/p_0_out [124]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[124]_i_1__0 
       (.I0(\r2/t0/t0/p_1_in [4]),
        .I1(\r2/t2/t2/p_0_in [4]),
        .I2(\r2/t1/t1/p_1_in [4]),
        .I3(\r2/t1/t1/p_0_in [4]),
        .I4(k1b[124]),
        .I5(\r2/t3/t3/p_0_in [4]),
        .O(\r2/p_0_out [124]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[124]_i_1__1 
       (.I0(\r3/t0/t0/p_1_in [4]),
        .I1(\r3/t2/t2/p_0_in [4]),
        .I2(\r3/t1/t1/p_1_in [4]),
        .I3(\r3/t1/t1/p_0_in [4]),
        .I4(k2b[124]),
        .I5(\r3/t3/t3/p_0_in [4]),
        .O(\r3/p_0_out [124]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[124]_i_1__2 
       (.I0(\r4/t0/t0/p_1_in [4]),
        .I1(\r4/t2/t2/p_0_in [4]),
        .I2(\r4/t1/t1/p_1_in [4]),
        .I3(\r4/t1/t1/p_0_in [4]),
        .I4(k3b[124]),
        .I5(\r4/t3/t3/p_0_in [4]),
        .O(\r4/p_0_out [124]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[124]_i_1__3 
       (.I0(\r5/t0/t0/p_1_in [4]),
        .I1(\r5/t2/t2/p_0_in [4]),
        .I2(\r5/t1/t1/p_1_in [4]),
        .I3(\r5/t1/t1/p_0_in [4]),
        .I4(k4b[124]),
        .I5(\r5/t3/t3/p_0_in [4]),
        .O(\r5/p_0_out [124]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[124]_i_1__4 
       (.I0(\r6/t0/t0/p_1_in [4]),
        .I1(\r6/t2/t2/p_0_in [4]),
        .I2(\r6/t1/t1/p_1_in [4]),
        .I3(\r6/t1/t1/p_0_in [4]),
        .I4(k5b[124]),
        .I5(\r6/t3/t3/p_0_in [4]),
        .O(\r6/p_0_out [124]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[124]_i_1__5 
       (.I0(\r7/t0/t0/p_1_in [4]),
        .I1(\r7/t2/t2/p_0_in [4]),
        .I2(\r7/t1/t1/p_1_in [4]),
        .I3(\r7/t1/t1/p_0_in [4]),
        .I4(k6b[124]),
        .I5(\r7/t3/t3/p_0_in [4]),
        .O(\r7/p_0_out [124]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[124]_i_1__6 
       (.I0(\r8/t0/t0/p_1_in [4]),
        .I1(\r8/t2/t2/p_0_in [4]),
        .I2(\r8/t1/t1/p_1_in [4]),
        .I3(\r8/t1/t1/p_0_in [4]),
        .I4(k7b[124]),
        .I5(\r8/t3/t3/p_0_in [4]),
        .O(\r8/p_0_out [124]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[124]_i_1__7 
       (.I0(\r9/t0/t0/p_1_in [4]),
        .I1(\r9/t2/t2/p_0_in [4]),
        .I2(\r9/t1/t1/p_1_in [4]),
        .I3(\r9/t1/t1/p_0_in [4]),
        .I4(k8b[124]),
        .I5(\r9/t3/t3/p_0_in [4]),
        .O(\r9/p_0_out [124]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair320" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[124]_i_1__8 
       (.I0(\a10/k0a [28]),
        .I1(\a10/k4a [28]),
        .I2(\rf/p_3_in [28]),
        .O(\rf/p_4_out [124]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[125]_i_1 
       (.I0(\r1/t0/t0/p_1_in [5]),
        .I1(\r1/t2/t2/p_0_in [5]),
        .I2(\r1/t1/t1/p_1_in [5]),
        .I3(\r1/t1/t1/p_0_in [5]),
        .I4(k0b[125]),
        .I5(\r1/t3/t3/p_0_in [5]),
        .O(\r1/p_0_out [125]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[125]_i_1__0 
       (.I0(\r2/t0/t0/p_1_in [5]),
        .I1(\r2/t2/t2/p_0_in [5]),
        .I2(\r2/t1/t1/p_1_in [5]),
        .I3(\r2/t1/t1/p_0_in [5]),
        .I4(k1b[125]),
        .I5(\r2/t3/t3/p_0_in [5]),
        .O(\r2/p_0_out [125]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[125]_i_1__1 
       (.I0(\r3/t0/t0/p_1_in [5]),
        .I1(\r3/t2/t2/p_0_in [5]),
        .I2(\r3/t1/t1/p_1_in [5]),
        .I3(\r3/t1/t1/p_0_in [5]),
        .I4(k2b[125]),
        .I5(\r3/t3/t3/p_0_in [5]),
        .O(\r3/p_0_out [125]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[125]_i_1__2 
       (.I0(\r4/t0/t0/p_1_in [5]),
        .I1(\r4/t2/t2/p_0_in [5]),
        .I2(\r4/t1/t1/p_1_in [5]),
        .I3(\r4/t1/t1/p_0_in [5]),
        .I4(k3b[125]),
        .I5(\r4/t3/t3/p_0_in [5]),
        .O(\r4/p_0_out [125]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[125]_i_1__3 
       (.I0(\r5/t0/t0/p_1_in [5]),
        .I1(\r5/t2/t2/p_0_in [5]),
        .I2(\r5/t1/t1/p_1_in [5]),
        .I3(\r5/t1/t1/p_0_in [5]),
        .I4(k4b[125]),
        .I5(\r5/t3/t3/p_0_in [5]),
        .O(\r5/p_0_out [125]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[125]_i_1__4 
       (.I0(\r6/t0/t0/p_1_in [5]),
        .I1(\r6/t2/t2/p_0_in [5]),
        .I2(\r6/t1/t1/p_1_in [5]),
        .I3(\r6/t1/t1/p_0_in [5]),
        .I4(k5b[125]),
        .I5(\r6/t3/t3/p_0_in [5]),
        .O(\r6/p_0_out [125]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[125]_i_1__5 
       (.I0(\r7/t0/t0/p_1_in [5]),
        .I1(\r7/t2/t2/p_0_in [5]),
        .I2(\r7/t1/t1/p_1_in [5]),
        .I3(\r7/t1/t1/p_0_in [5]),
        .I4(k6b[125]),
        .I5(\r7/t3/t3/p_0_in [5]),
        .O(\r7/p_0_out [125]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[125]_i_1__6 
       (.I0(\r8/t0/t0/p_1_in [5]),
        .I1(\r8/t2/t2/p_0_in [5]),
        .I2(\r8/t1/t1/p_1_in [5]),
        .I3(\r8/t1/t1/p_0_in [5]),
        .I4(k7b[125]),
        .I5(\r8/t3/t3/p_0_in [5]),
        .O(\r8/p_0_out [125]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[125]_i_1__7 
       (.I0(\r9/t0/t0/p_1_in [5]),
        .I1(\r9/t2/t2/p_0_in [5]),
        .I2(\r9/t1/t1/p_1_in [5]),
        .I3(\r9/t1/t1/p_0_in [5]),
        .I4(k8b[125]),
        .I5(\r9/t3/t3/p_0_in [5]),
        .O(\r9/p_0_out [125]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair321" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[125]_i_1__8 
       (.I0(\a10/k0a [29]),
        .I1(\a10/k4a [29]),
        .I2(\rf/p_3_in [29]),
        .O(\rf/p_4_out [125]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[126]_i_1 
       (.I0(\r1/t0/t0/p_1_in [6]),
        .I1(\r1/t2/t2/p_0_in [6]),
        .I2(\r1/t1/t1/p_1_in [6]),
        .I3(\r1/t1/t1/p_0_in [6]),
        .I4(k0b[126]),
        .I5(\r1/t3/t3/p_0_in [6]),
        .O(\r1/p_0_out [126]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[126]_i_1__0 
       (.I0(\r2/t0/t0/p_1_in [6]),
        .I1(\r2/t2/t2/p_0_in [6]),
        .I2(\r2/t1/t1/p_1_in [6]),
        .I3(\r2/t1/t1/p_0_in [6]),
        .I4(k1b[126]),
        .I5(\r2/t3/t3/p_0_in [6]),
        .O(\r2/p_0_out [126]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[126]_i_1__1 
       (.I0(\r3/t0/t0/p_1_in [6]),
        .I1(\r3/t2/t2/p_0_in [6]),
        .I2(\r3/t1/t1/p_1_in [6]),
        .I3(\r3/t1/t1/p_0_in [6]),
        .I4(k2b[126]),
        .I5(\r3/t3/t3/p_0_in [6]),
        .O(\r3/p_0_out [126]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[126]_i_1__2 
       (.I0(\r4/t0/t0/p_1_in [6]),
        .I1(\r4/t2/t2/p_0_in [6]),
        .I2(\r4/t1/t1/p_1_in [6]),
        .I3(\r4/t1/t1/p_0_in [6]),
        .I4(k3b[126]),
        .I5(\r4/t3/t3/p_0_in [6]),
        .O(\r4/p_0_out [126]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[126]_i_1__3 
       (.I0(\r5/t0/t0/p_1_in [6]),
        .I1(\r5/t2/t2/p_0_in [6]),
        .I2(\r5/t1/t1/p_1_in [6]),
        .I3(\r5/t1/t1/p_0_in [6]),
        .I4(k4b[126]),
        .I5(\r5/t3/t3/p_0_in [6]),
        .O(\r5/p_0_out [126]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[126]_i_1__4 
       (.I0(\r6/t0/t0/p_1_in [6]),
        .I1(\r6/t2/t2/p_0_in [6]),
        .I2(\r6/t1/t1/p_1_in [6]),
        .I3(\r6/t1/t1/p_0_in [6]),
        .I4(k5b[126]),
        .I5(\r6/t3/t3/p_0_in [6]),
        .O(\r6/p_0_out [126]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[126]_i_1__5 
       (.I0(\r7/t0/t0/p_1_in [6]),
        .I1(\r7/t2/t2/p_0_in [6]),
        .I2(\r7/t1/t1/p_1_in [6]),
        .I3(\r7/t1/t1/p_0_in [6]),
        .I4(k6b[126]),
        .I5(\r7/t3/t3/p_0_in [6]),
        .O(\r7/p_0_out [126]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[126]_i_1__6 
       (.I0(\r8/t0/t0/p_1_in [6]),
        .I1(\r8/t2/t2/p_0_in [6]),
        .I2(\r8/t1/t1/p_1_in [6]),
        .I3(\r8/t1/t1/p_0_in [6]),
        .I4(k7b[126]),
        .I5(\r8/t3/t3/p_0_in [6]),
        .O(\r8/p_0_out [126]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[126]_i_1__7 
       (.I0(\r9/t0/t0/p_1_in [6]),
        .I1(\r9/t2/t2/p_0_in [6]),
        .I2(\r9/t1/t1/p_1_in [6]),
        .I3(\r9/t1/t1/p_0_in [6]),
        .I4(k8b[126]),
        .I5(\r9/t3/t3/p_0_in [6]),
        .O(\r9/p_0_out [126]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair323" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[126]_i_1__8 
       (.I0(\a10/k0a [30]),
        .I1(\a10/k4a [30]),
        .I2(\rf/p_3_in [30]),
        .O(\rf/p_4_out [126]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[127]_i_1 
       (.I0(\r1/t0/t0/p_1_in [7]),
        .I1(\r1/t2/t2/p_0_in [7]),
        .I2(\r1/t1/t1/p_1_in [7]),
        .I3(\r1/t1/t1/p_0_in [7]),
        .I4(k0b[127]),
        .I5(\r1/t3/t3/p_0_in [7]),
        .O(\r1/p_0_out [127]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[127]_i_1__0 
       (.I0(\r2/t0/t0/p_1_in [7]),
        .I1(\r2/t2/t2/p_0_in [7]),
        .I2(\r2/t1/t1/p_1_in [7]),
        .I3(\r2/t1/t1/p_0_in [7]),
        .I4(k1b[127]),
        .I5(\r2/t3/t3/p_0_in [7]),
        .O(\r2/p_0_out [127]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[127]_i_1__1 
       (.I0(\r3/t0/t0/p_1_in [7]),
        .I1(\r3/t2/t2/p_0_in [7]),
        .I2(\r3/t1/t1/p_1_in [7]),
        .I3(\r3/t1/t1/p_0_in [7]),
        .I4(k2b[127]),
        .I5(\r3/t3/t3/p_0_in [7]),
        .O(\r3/p_0_out [127]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[127]_i_1__2 
       (.I0(\r4/t0/t0/p_1_in [7]),
        .I1(\r4/t2/t2/p_0_in [7]),
        .I2(\r4/t1/t1/p_1_in [7]),
        .I3(\r4/t1/t1/p_0_in [7]),
        .I4(k3b[127]),
        .I5(\r4/t3/t3/p_0_in [7]),
        .O(\r4/p_0_out [127]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[127]_i_1__3 
       (.I0(\r5/t0/t0/p_1_in [7]),
        .I1(\r5/t2/t2/p_0_in [7]),
        .I2(\r5/t1/t1/p_1_in [7]),
        .I3(\r5/t1/t1/p_0_in [7]),
        .I4(k4b[127]),
        .I5(\r5/t3/t3/p_0_in [7]),
        .O(\r5/p_0_out [127]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[127]_i_1__4 
       (.I0(\r6/t0/t0/p_1_in [7]),
        .I1(\r6/t2/t2/p_0_in [7]),
        .I2(\r6/t1/t1/p_1_in [7]),
        .I3(\r6/t1/t1/p_0_in [7]),
        .I4(k5b[127]),
        .I5(\r6/t3/t3/p_0_in [7]),
        .O(\r6/p_0_out [127]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[127]_i_1__5 
       (.I0(\r7/t0/t0/p_1_in [7]),
        .I1(\r7/t2/t2/p_0_in [7]),
        .I2(\r7/t1/t1/p_1_in [7]),
        .I3(\r7/t1/t1/p_0_in [7]),
        .I4(k6b[127]),
        .I5(\r7/t3/t3/p_0_in [7]),
        .O(\r7/p_0_out [127]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[127]_i_1__6 
       (.I0(\r8/t0/t0/p_1_in [7]),
        .I1(\r8/t2/t2/p_0_in [7]),
        .I2(\r8/t1/t1/p_1_in [7]),
        .I3(\r8/t1/t1/p_0_in [7]),
        .I4(k7b[127]),
        .I5(\r8/t3/t3/p_0_in [7]),
        .O(\r8/p_0_out [127]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[127]_i_1__7 
       (.I0(\r9/t0/t0/p_1_in [7]),
        .I1(\r9/t2/t2/p_0_in [7]),
        .I2(\r9/t1/t1/p_1_in [7]),
        .I3(\r9/t1/t1/p_0_in [7]),
        .I4(k8b[127]),
        .I5(\r9/t3/t3/p_0_in [7]),
        .O(\r9/p_0_out [127]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair324" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[127]_i_1__8 
       (.I0(\a10/k0a [31]),
        .I1(\a10/k4a [31]),
        .I2(\rf/p_3_in [31]),
        .O(\rf/p_4_out [127]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[12]_i_1 
       (.I0(\r1/t0/t1/p_0_in [4]),
        .I1(\r1/t2/t3/p_1_in [4]),
        .I2(\r1/t2/t3/p_0_in [4]),
        .I3(\r1/t1/t2/p_1_in [4]),
        .I4(k0b[12]),
        .I5(\r1/t3/t0/p_0_in [4]),
        .O(\r1/p_0_out [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[12]_i_1__0 
       (.I0(\r2/t0/t1/p_0_in [4]),
        .I1(\r2/t2/t3/p_1_in [4]),
        .I2(\r2/t2/t3/p_0_in [4]),
        .I3(\r2/t1/t2/p_1_in [4]),
        .I4(k1b[12]),
        .I5(\r2/t3/t0/p_0_in [4]),
        .O(\r2/p_0_out [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[12]_i_1__1 
       (.I0(\r3/t0/t1/p_0_in [4]),
        .I1(\r3/t2/t3/p_1_in [4]),
        .I2(\r3/t2/t3/p_0_in [4]),
        .I3(\r3/t1/t2/p_1_in [4]),
        .I4(k2b[12]),
        .I5(\r3/t3/t0/p_0_in [4]),
        .O(\r3/p_0_out [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[12]_i_1__2 
       (.I0(\r4/t0/t1/p_0_in [4]),
        .I1(\r4/t2/t3/p_1_in [4]),
        .I2(\r4/t2/t3/p_0_in [4]),
        .I3(\r4/t1/t2/p_1_in [4]),
        .I4(k3b[12]),
        .I5(\r4/t3/t0/p_0_in [4]),
        .O(\r4/p_0_out [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[12]_i_1__3 
       (.I0(\r5/t0/t1/p_0_in [4]),
        .I1(\r5/t2/t3/p_1_in [4]),
        .I2(\r5/t2/t3/p_0_in [4]),
        .I3(\r5/t1/t2/p_1_in [4]),
        .I4(k4b[12]),
        .I5(\r5/t3/t0/p_0_in [4]),
        .O(\r5/p_0_out [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[12]_i_1__4 
       (.I0(\r6/t0/t1/p_0_in [4]),
        .I1(\r6/t2/t3/p_1_in [4]),
        .I2(\r6/t2/t3/p_0_in [4]),
        .I3(\r6/t1/t2/p_1_in [4]),
        .I4(k5b[12]),
        .I5(\r6/t3/t0/p_0_in [4]),
        .O(\r6/p_0_out [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[12]_i_1__5 
       (.I0(\r7/t0/t1/p_0_in [4]),
        .I1(\r7/t2/t3/p_1_in [4]),
        .I2(\r7/t2/t3/p_0_in [4]),
        .I3(\r7/t1/t2/p_1_in [4]),
        .I4(k6b[12]),
        .I5(\r7/t3/t0/p_0_in [4]),
        .O(\r7/p_0_out [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[12]_i_1__6 
       (.I0(\r8/t0/t1/p_0_in [4]),
        .I1(\r8/t2/t3/p_1_in [4]),
        .I2(\r8/t2/t3/p_0_in [4]),
        .I3(\r8/t1/t2/p_1_in [4]),
        .I4(k7b[12]),
        .I5(\r8/t3/t0/p_0_in [4]),
        .O(\r8/p_0_out [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[12]_i_1__7 
       (.I0(\r9/t0/t1/p_0_in [4]),
        .I1(\r9/t2/t3/p_1_in [4]),
        .I2(\r9/t2/t3/p_0_in [4]),
        .I3(\r9/t1/t2/p_1_in [4]),
        .I4(k8b[12]),
        .I5(\r9/t3/t0/p_0_in [4]),
        .O(\r9/p_0_out [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair330" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[12]_i_1__8 
       (.I0(\a10/k3a [12]),
        .I1(\a10/k4a [12]),
        .I2(\rf/p_0_in [12]),
        .O(\rf/p_4_out [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[13]_i_1 
       (.I0(\r1/t0/t1/p_0_in [5]),
        .I1(\r1/t2/t3/p_1_in [5]),
        .I2(\r1/t2/t3/p_0_in [5]),
        .I3(\r1/t1/t2/p_1_in [5]),
        .I4(k0b[13]),
        .I5(\r1/t3/t0/p_0_in [5]),
        .O(\r1/p_0_out [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[13]_i_1__0 
       (.I0(\r2/t0/t1/p_0_in [5]),
        .I1(\r2/t2/t3/p_1_in [5]),
        .I2(\r2/t2/t3/p_0_in [5]),
        .I3(\r2/t1/t2/p_1_in [5]),
        .I4(k1b[13]),
        .I5(\r2/t3/t0/p_0_in [5]),
        .O(\r2/p_0_out [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[13]_i_1__1 
       (.I0(\r3/t0/t1/p_0_in [5]),
        .I1(\r3/t2/t3/p_1_in [5]),
        .I2(\r3/t2/t3/p_0_in [5]),
        .I3(\r3/t1/t2/p_1_in [5]),
        .I4(k2b[13]),
        .I5(\r3/t3/t0/p_0_in [5]),
        .O(\r3/p_0_out [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[13]_i_1__2 
       (.I0(\r4/t0/t1/p_0_in [5]),
        .I1(\r4/t2/t3/p_1_in [5]),
        .I2(\r4/t2/t3/p_0_in [5]),
        .I3(\r4/t1/t2/p_1_in [5]),
        .I4(k3b[13]),
        .I5(\r4/t3/t0/p_0_in [5]),
        .O(\r4/p_0_out [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[13]_i_1__3 
       (.I0(\r5/t0/t1/p_0_in [5]),
        .I1(\r5/t2/t3/p_1_in [5]),
        .I2(\r5/t2/t3/p_0_in [5]),
        .I3(\r5/t1/t2/p_1_in [5]),
        .I4(k4b[13]),
        .I5(\r5/t3/t0/p_0_in [5]),
        .O(\r5/p_0_out [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[13]_i_1__4 
       (.I0(\r6/t0/t1/p_0_in [5]),
        .I1(\r6/t2/t3/p_1_in [5]),
        .I2(\r6/t2/t3/p_0_in [5]),
        .I3(\r6/t1/t2/p_1_in [5]),
        .I4(k5b[13]),
        .I5(\r6/t3/t0/p_0_in [5]),
        .O(\r6/p_0_out [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[13]_i_1__5 
       (.I0(\r7/t0/t1/p_0_in [5]),
        .I1(\r7/t2/t3/p_1_in [5]),
        .I2(\r7/t2/t3/p_0_in [5]),
        .I3(\r7/t1/t2/p_1_in [5]),
        .I4(k6b[13]),
        .I5(\r7/t3/t0/p_0_in [5]),
        .O(\r7/p_0_out [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[13]_i_1__6 
       (.I0(\r8/t0/t1/p_0_in [5]),
        .I1(\r8/t2/t3/p_1_in [5]),
        .I2(\r8/t2/t3/p_0_in [5]),
        .I3(\r8/t1/t2/p_1_in [5]),
        .I4(k7b[13]),
        .I5(\r8/t3/t0/p_0_in [5]),
        .O(\r8/p_0_out [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[13]_i_1__7 
       (.I0(\r9/t0/t1/p_0_in [5]),
        .I1(\r9/t2/t3/p_1_in [5]),
        .I2(\r9/t2/t3/p_0_in [5]),
        .I3(\r9/t1/t2/p_1_in [5]),
        .I4(k8b[13]),
        .I5(\r9/t3/t0/p_0_in [5]),
        .O(\r9/p_0_out [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair329" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[13]_i_1__8 
       (.I0(\a10/k3a [13]),
        .I1(\a10/k4a [13]),
        .I2(\rf/p_0_in [13]),
        .O(\rf/p_4_out [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[14]_i_1 
       (.I0(\r1/t0/t1/p_0_in [6]),
        .I1(\r1/t2/t3/p_1_in [6]),
        .I2(\r1/t2/t3/p_0_in [6]),
        .I3(\r1/t1/t2/p_1_in [6]),
        .I4(k0b[14]),
        .I5(\r1/t3/t0/p_0_in [6]),
        .O(\r1/p_0_out [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[14]_i_1__0 
       (.I0(\r2/t0/t1/p_0_in [6]),
        .I1(\r2/t2/t3/p_1_in [6]),
        .I2(\r2/t2/t3/p_0_in [6]),
        .I3(\r2/t1/t2/p_1_in [6]),
        .I4(k1b[14]),
        .I5(\r2/t3/t0/p_0_in [6]),
        .O(\r2/p_0_out [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[14]_i_1__1 
       (.I0(\r3/t0/t1/p_0_in [6]),
        .I1(\r3/t2/t3/p_1_in [6]),
        .I2(\r3/t2/t3/p_0_in [6]),
        .I3(\r3/t1/t2/p_1_in [6]),
        .I4(k2b[14]),
        .I5(\r3/t3/t0/p_0_in [6]),
        .O(\r3/p_0_out [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[14]_i_1__2 
       (.I0(\r4/t0/t1/p_0_in [6]),
        .I1(\r4/t2/t3/p_1_in [6]),
        .I2(\r4/t2/t3/p_0_in [6]),
        .I3(\r4/t1/t2/p_1_in [6]),
        .I4(k3b[14]),
        .I5(\r4/t3/t0/p_0_in [6]),
        .O(\r4/p_0_out [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[14]_i_1__3 
       (.I0(\r5/t0/t1/p_0_in [6]),
        .I1(\r5/t2/t3/p_1_in [6]),
        .I2(\r5/t2/t3/p_0_in [6]),
        .I3(\r5/t1/t2/p_1_in [6]),
        .I4(k4b[14]),
        .I5(\r5/t3/t0/p_0_in [6]),
        .O(\r5/p_0_out [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[14]_i_1__4 
       (.I0(\r6/t0/t1/p_0_in [6]),
        .I1(\r6/t2/t3/p_1_in [6]),
        .I2(\r6/t2/t3/p_0_in [6]),
        .I3(\r6/t1/t2/p_1_in [6]),
        .I4(k5b[14]),
        .I5(\r6/t3/t0/p_0_in [6]),
        .O(\r6/p_0_out [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[14]_i_1__5 
       (.I0(\r7/t0/t1/p_0_in [6]),
        .I1(\r7/t2/t3/p_1_in [6]),
        .I2(\r7/t2/t3/p_0_in [6]),
        .I3(\r7/t1/t2/p_1_in [6]),
        .I4(k6b[14]),
        .I5(\r7/t3/t0/p_0_in [6]),
        .O(\r7/p_0_out [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[14]_i_1__6 
       (.I0(\r8/t0/t1/p_0_in [6]),
        .I1(\r8/t2/t3/p_1_in [6]),
        .I2(\r8/t2/t3/p_0_in [6]),
        .I3(\r8/t1/t2/p_1_in [6]),
        .I4(k7b[14]),
        .I5(\r8/t3/t0/p_0_in [6]),
        .O(\r8/p_0_out [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[14]_i_1__7 
       (.I0(\r9/t0/t1/p_0_in [6]),
        .I1(\r9/t2/t3/p_1_in [6]),
        .I2(\r9/t2/t3/p_0_in [6]),
        .I3(\r9/t1/t2/p_1_in [6]),
        .I4(k8b[14]),
        .I5(\r9/t3/t0/p_0_in [6]),
        .O(\r9/p_0_out [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair328" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[14]_i_1__8 
       (.I0(\a10/k3a [14]),
        .I1(\a10/k4a [14]),
        .I2(\rf/p_0_in [14]),
        .O(\rf/p_4_out [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[15]_i_1 
       (.I0(\r1/t0/t1/p_0_in [7]),
        .I1(\r1/t2/t3/p_1_in [7]),
        .I2(\r1/t2/t3/p_0_in [7]),
        .I3(\r1/t1/t2/p_1_in [7]),
        .I4(k0b[15]),
        .I5(\r1/t3/t0/p_0_in [7]),
        .O(\r1/p_0_out [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[15]_i_1__0 
       (.I0(\r2/t0/t1/p_0_in [7]),
        .I1(\r2/t2/t3/p_1_in [7]),
        .I2(\r2/t2/t3/p_0_in [7]),
        .I3(\r2/t1/t2/p_1_in [7]),
        .I4(k1b[15]),
        .I5(\r2/t3/t0/p_0_in [7]),
        .O(\r2/p_0_out [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[15]_i_1__1 
       (.I0(\r3/t0/t1/p_0_in [7]),
        .I1(\r3/t2/t3/p_1_in [7]),
        .I2(\r3/t2/t3/p_0_in [7]),
        .I3(\r3/t1/t2/p_1_in [7]),
        .I4(k2b[15]),
        .I5(\r3/t3/t0/p_0_in [7]),
        .O(\r3/p_0_out [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[15]_i_1__2 
       (.I0(\r4/t0/t1/p_0_in [7]),
        .I1(\r4/t2/t3/p_1_in [7]),
        .I2(\r4/t2/t3/p_0_in [7]),
        .I3(\r4/t1/t2/p_1_in [7]),
        .I4(k3b[15]),
        .I5(\r4/t3/t0/p_0_in [7]),
        .O(\r4/p_0_out [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[15]_i_1__3 
       (.I0(\r5/t0/t1/p_0_in [7]),
        .I1(\r5/t2/t3/p_1_in [7]),
        .I2(\r5/t2/t3/p_0_in [7]),
        .I3(\r5/t1/t2/p_1_in [7]),
        .I4(k4b[15]),
        .I5(\r5/t3/t0/p_0_in [7]),
        .O(\r5/p_0_out [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[15]_i_1__4 
       (.I0(\r6/t0/t1/p_0_in [7]),
        .I1(\r6/t2/t3/p_1_in [7]),
        .I2(\r6/t2/t3/p_0_in [7]),
        .I3(\r6/t1/t2/p_1_in [7]),
        .I4(k5b[15]),
        .I5(\r6/t3/t0/p_0_in [7]),
        .O(\r6/p_0_out [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[15]_i_1__5 
       (.I0(\r7/t0/t1/p_0_in [7]),
        .I1(\r7/t2/t3/p_1_in [7]),
        .I2(\r7/t2/t3/p_0_in [7]),
        .I3(\r7/t1/t2/p_1_in [7]),
        .I4(k6b[15]),
        .I5(\r7/t3/t0/p_0_in [7]),
        .O(\r7/p_0_out [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[15]_i_1__6 
       (.I0(\r8/t0/t1/p_0_in [7]),
        .I1(\r8/t2/t3/p_1_in [7]),
        .I2(\r8/t2/t3/p_0_in [7]),
        .I3(\r8/t1/t2/p_1_in [7]),
        .I4(k7b[15]),
        .I5(\r8/t3/t0/p_0_in [7]),
        .O(\r8/p_0_out [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[15]_i_1__7 
       (.I0(\r9/t0/t1/p_0_in [7]),
        .I1(\r9/t2/t3/p_1_in [7]),
        .I2(\r9/t2/t3/p_0_in [7]),
        .I3(\r9/t1/t2/p_1_in [7]),
        .I4(k8b[15]),
        .I5(\r9/t3/t0/p_0_in [7]),
        .O(\r9/p_0_out [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair359" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[15]_i_1__8 
       (.I0(\a10/k3a [15]),
        .I1(\a10/k4a [15]),
        .I2(\rf/p_0_in [15]),
        .O(\rf/p_4_out [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[16]_i_1 
       (.I0(\r1/t0/t1/p_1_in [0]),
        .I1(\r1/t2/t3/p_0_in [0]),
        .I2(\r1/t1/t2/p_1_in [0]),
        .I3(\r1/t1/t2/p_0_in [0]),
        .I4(k0b[16]),
        .I5(\r1/t3/t0/p_0_in [0]),
        .O(\r1/p_0_out [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[16]_i_1__0 
       (.I0(\r2/t0/t1/p_1_in [0]),
        .I1(\r2/t2/t3/p_0_in [0]),
        .I2(\r2/t1/t2/p_1_in [0]),
        .I3(\r2/t1/t2/p_0_in [0]),
        .I4(k1b[16]),
        .I5(\r2/t3/t0/p_0_in [0]),
        .O(\r2/p_0_out [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[16]_i_1__1 
       (.I0(\r3/t0/t1/p_1_in [0]),
        .I1(\r3/t2/t3/p_0_in [0]),
        .I2(\r3/t1/t2/p_1_in [0]),
        .I3(\r3/t1/t2/p_0_in [0]),
        .I4(k2b[16]),
        .I5(\r3/t3/t0/p_0_in [0]),
        .O(\r3/p_0_out [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[16]_i_1__2 
       (.I0(\r4/t0/t1/p_1_in [0]),
        .I1(\r4/t2/t3/p_0_in [0]),
        .I2(\r4/t1/t2/p_1_in [0]),
        .I3(\r4/t1/t2/p_0_in [0]),
        .I4(k3b[16]),
        .I5(\r4/t3/t0/p_0_in [0]),
        .O(\r4/p_0_out [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[16]_i_1__3 
       (.I0(\r5/t0/t1/p_1_in [0]),
        .I1(\r5/t2/t3/p_0_in [0]),
        .I2(\r5/t1/t2/p_1_in [0]),
        .I3(\r5/t1/t2/p_0_in [0]),
        .I4(k4b[16]),
        .I5(\r5/t3/t0/p_0_in [0]),
        .O(\r5/p_0_out [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[16]_i_1__4 
       (.I0(\r6/t0/t1/p_1_in [0]),
        .I1(\r6/t2/t3/p_0_in [0]),
        .I2(\r6/t1/t2/p_1_in [0]),
        .I3(\r6/t1/t2/p_0_in [0]),
        .I4(k5b[16]),
        .I5(\r6/t3/t0/p_0_in [0]),
        .O(\r6/p_0_out [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[16]_i_1__5 
       (.I0(\r7/t0/t1/p_1_in [0]),
        .I1(\r7/t2/t3/p_0_in [0]),
        .I2(\r7/t1/t2/p_1_in [0]),
        .I3(\r7/t1/t2/p_0_in [0]),
        .I4(k6b[16]),
        .I5(\r7/t3/t0/p_0_in [0]),
        .O(\r7/p_0_out [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[16]_i_1__6 
       (.I0(\r8/t0/t1/p_1_in [0]),
        .I1(\r8/t2/t3/p_0_in [0]),
        .I2(\r8/t1/t2/p_1_in [0]),
        .I3(\r8/t1/t2/p_0_in [0]),
        .I4(k7b[16]),
        .I5(\r8/t3/t0/p_0_in [0]),
        .O(\r8/p_0_out [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[16]_i_1__7 
       (.I0(\r9/t0/t1/p_1_in [0]),
        .I1(\r9/t2/t3/p_0_in [0]),
        .I2(\r9/t1/t2/p_1_in [0]),
        .I3(\r9/t1/t2/p_0_in [0]),
        .I4(k8b[16]),
        .I5(\r9/t3/t0/p_0_in [0]),
        .O(\r9/p_0_out [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair358" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[16]_i_1__8 
       (.I0(\a10/k3a [16]),
        .I1(\a10/k4a [16]),
        .I2(\rf/p_0_in [16]),
        .O(\rf/p_4_out [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[17]_i_1 
       (.I0(\r1/t0/t1/p_1_in [1]),
        .I1(\r1/t2/t3/p_0_in [1]),
        .I2(\r1/t1/t2/p_1_in [1]),
        .I3(\r1/t1/t2/p_0_in [1]),
        .I4(k0b[17]),
        .I5(\r1/t3/t0/p_0_in [1]),
        .O(\r1/p_0_out [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[17]_i_1__0 
       (.I0(\r2/t0/t1/p_1_in [1]),
        .I1(\r2/t2/t3/p_0_in [1]),
        .I2(\r2/t1/t2/p_1_in [1]),
        .I3(\r2/t1/t2/p_0_in [1]),
        .I4(k1b[17]),
        .I5(\r2/t3/t0/p_0_in [1]),
        .O(\r2/p_0_out [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[17]_i_1__1 
       (.I0(\r3/t0/t1/p_1_in [1]),
        .I1(\r3/t2/t3/p_0_in [1]),
        .I2(\r3/t1/t2/p_1_in [1]),
        .I3(\r3/t1/t2/p_0_in [1]),
        .I4(k2b[17]),
        .I5(\r3/t3/t0/p_0_in [1]),
        .O(\r3/p_0_out [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[17]_i_1__2 
       (.I0(\r4/t0/t1/p_1_in [1]),
        .I1(\r4/t2/t3/p_0_in [1]),
        .I2(\r4/t1/t2/p_1_in [1]),
        .I3(\r4/t1/t2/p_0_in [1]),
        .I4(k3b[17]),
        .I5(\r4/t3/t0/p_0_in [1]),
        .O(\r4/p_0_out [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[17]_i_1__3 
       (.I0(\r5/t0/t1/p_1_in [1]),
        .I1(\r5/t2/t3/p_0_in [1]),
        .I2(\r5/t1/t2/p_1_in [1]),
        .I3(\r5/t1/t2/p_0_in [1]),
        .I4(k4b[17]),
        .I5(\r5/t3/t0/p_0_in [1]),
        .O(\r5/p_0_out [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[17]_i_1__4 
       (.I0(\r6/t0/t1/p_1_in [1]),
        .I1(\r6/t2/t3/p_0_in [1]),
        .I2(\r6/t1/t2/p_1_in [1]),
        .I3(\r6/t1/t2/p_0_in [1]),
        .I4(k5b[17]),
        .I5(\r6/t3/t0/p_0_in [1]),
        .O(\r6/p_0_out [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[17]_i_1__5 
       (.I0(\r7/t0/t1/p_1_in [1]),
        .I1(\r7/t2/t3/p_0_in [1]),
        .I2(\r7/t1/t2/p_1_in [1]),
        .I3(\r7/t1/t2/p_0_in [1]),
        .I4(k6b[17]),
        .I5(\r7/t3/t0/p_0_in [1]),
        .O(\r7/p_0_out [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[17]_i_1__6 
       (.I0(\r8/t0/t1/p_1_in [1]),
        .I1(\r8/t2/t3/p_0_in [1]),
        .I2(\r8/t1/t2/p_1_in [1]),
        .I3(\r8/t1/t2/p_0_in [1]),
        .I4(k7b[17]),
        .I5(\r8/t3/t0/p_0_in [1]),
        .O(\r8/p_0_out [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[17]_i_1__7 
       (.I0(\r9/t0/t1/p_1_in [1]),
        .I1(\r9/t2/t3/p_0_in [1]),
        .I2(\r9/t1/t2/p_1_in [1]),
        .I3(\r9/t1/t2/p_0_in [1]),
        .I4(k8b[17]),
        .I5(\r9/t3/t0/p_0_in [1]),
        .O(\r9/p_0_out [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair357" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[17]_i_1__8 
       (.I0(\a10/k3a [17]),
        .I1(\a10/k4a [17]),
        .I2(\rf/p_0_in [17]),
        .O(\rf/p_4_out [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[18]_i_1 
       (.I0(\r1/t0/t1/p_1_in [2]),
        .I1(\r1/t2/t3/p_0_in [2]),
        .I2(\r1/t1/t2/p_1_in [2]),
        .I3(\r1/t1/t2/p_0_in [2]),
        .I4(k0b[18]),
        .I5(\r1/t3/t0/p_0_in [2]),
        .O(\r1/p_0_out [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[18]_i_1__0 
       (.I0(\r2/t0/t1/p_1_in [2]),
        .I1(\r2/t2/t3/p_0_in [2]),
        .I2(\r2/t1/t2/p_1_in [2]),
        .I3(\r2/t1/t2/p_0_in [2]),
        .I4(k1b[18]),
        .I5(\r2/t3/t0/p_0_in [2]),
        .O(\r2/p_0_out [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[18]_i_1__1 
       (.I0(\r3/t0/t1/p_1_in [2]),
        .I1(\r3/t2/t3/p_0_in [2]),
        .I2(\r3/t1/t2/p_1_in [2]),
        .I3(\r3/t1/t2/p_0_in [2]),
        .I4(k2b[18]),
        .I5(\r3/t3/t0/p_0_in [2]),
        .O(\r3/p_0_out [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[18]_i_1__2 
       (.I0(\r4/t0/t1/p_1_in [2]),
        .I1(\r4/t2/t3/p_0_in [2]),
        .I2(\r4/t1/t2/p_1_in [2]),
        .I3(\r4/t1/t2/p_0_in [2]),
        .I4(k3b[18]),
        .I5(\r4/t3/t0/p_0_in [2]),
        .O(\r4/p_0_out [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[18]_i_1__3 
       (.I0(\r5/t0/t1/p_1_in [2]),
        .I1(\r5/t2/t3/p_0_in [2]),
        .I2(\r5/t1/t2/p_1_in [2]),
        .I3(\r5/t1/t2/p_0_in [2]),
        .I4(k4b[18]),
        .I5(\r5/t3/t0/p_0_in [2]),
        .O(\r5/p_0_out [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[18]_i_1__4 
       (.I0(\r6/t0/t1/p_1_in [2]),
        .I1(\r6/t2/t3/p_0_in [2]),
        .I2(\r6/t1/t2/p_1_in [2]),
        .I3(\r6/t1/t2/p_0_in [2]),
        .I4(k5b[18]),
        .I5(\r6/t3/t0/p_0_in [2]),
        .O(\r6/p_0_out [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[18]_i_1__5 
       (.I0(\r7/t0/t1/p_1_in [2]),
        .I1(\r7/t2/t3/p_0_in [2]),
        .I2(\r7/t1/t2/p_1_in [2]),
        .I3(\r7/t1/t2/p_0_in [2]),
        .I4(k6b[18]),
        .I5(\r7/t3/t0/p_0_in [2]),
        .O(\r7/p_0_out [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[18]_i_1__6 
       (.I0(\r8/t0/t1/p_1_in [2]),
        .I1(\r8/t2/t3/p_0_in [2]),
        .I2(\r8/t1/t2/p_1_in [2]),
        .I3(\r8/t1/t2/p_0_in [2]),
        .I4(k7b[18]),
        .I5(\r8/t3/t0/p_0_in [2]),
        .O(\r8/p_0_out [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[18]_i_1__7 
       (.I0(\r9/t0/t1/p_1_in [2]),
        .I1(\r9/t2/t3/p_0_in [2]),
        .I2(\r9/t1/t2/p_1_in [2]),
        .I3(\r9/t1/t2/p_0_in [2]),
        .I4(k8b[18]),
        .I5(\r9/t3/t0/p_0_in [2]),
        .O(\r9/p_0_out [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair356" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[18]_i_1__8 
       (.I0(\a10/k3a [18]),
        .I1(\a10/k4a [18]),
        .I2(\rf/p_0_in [18]),
        .O(\rf/p_4_out [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[19]_i_1 
       (.I0(\r1/t0/t1/p_1_in [3]),
        .I1(\r1/t2/t3/p_0_in [3]),
        .I2(\r1/t1/t2/p_1_in [3]),
        .I3(\r1/t1/t2/p_0_in [3]),
        .I4(k0b[19]),
        .I5(\r1/t3/t0/p_0_in [3]),
        .O(\r1/p_0_out [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[19]_i_1__0 
       (.I0(\r2/t0/t1/p_1_in [3]),
        .I1(\r2/t2/t3/p_0_in [3]),
        .I2(\r2/t1/t2/p_1_in [3]),
        .I3(\r2/t1/t2/p_0_in [3]),
        .I4(k1b[19]),
        .I5(\r2/t3/t0/p_0_in [3]),
        .O(\r2/p_0_out [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[19]_i_1__1 
       (.I0(\r3/t0/t1/p_1_in [3]),
        .I1(\r3/t2/t3/p_0_in [3]),
        .I2(\r3/t1/t2/p_1_in [3]),
        .I3(\r3/t1/t2/p_0_in [3]),
        .I4(k2b[19]),
        .I5(\r3/t3/t0/p_0_in [3]),
        .O(\r3/p_0_out [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[19]_i_1__2 
       (.I0(\r4/t0/t1/p_1_in [3]),
        .I1(\r4/t2/t3/p_0_in [3]),
        .I2(\r4/t1/t2/p_1_in [3]),
        .I3(\r4/t1/t2/p_0_in [3]),
        .I4(k3b[19]),
        .I5(\r4/t3/t0/p_0_in [3]),
        .O(\r4/p_0_out [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[19]_i_1__3 
       (.I0(\r5/t0/t1/p_1_in [3]),
        .I1(\r5/t2/t3/p_0_in [3]),
        .I2(\r5/t1/t2/p_1_in [3]),
        .I3(\r5/t1/t2/p_0_in [3]),
        .I4(k4b[19]),
        .I5(\r5/t3/t0/p_0_in [3]),
        .O(\r5/p_0_out [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[19]_i_1__4 
       (.I0(\r6/t0/t1/p_1_in [3]),
        .I1(\r6/t2/t3/p_0_in [3]),
        .I2(\r6/t1/t2/p_1_in [3]),
        .I3(\r6/t1/t2/p_0_in [3]),
        .I4(k5b[19]),
        .I5(\r6/t3/t0/p_0_in [3]),
        .O(\r6/p_0_out [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[19]_i_1__5 
       (.I0(\r7/t0/t1/p_1_in [3]),
        .I1(\r7/t2/t3/p_0_in [3]),
        .I2(\r7/t1/t2/p_1_in [3]),
        .I3(\r7/t1/t2/p_0_in [3]),
        .I4(k6b[19]),
        .I5(\r7/t3/t0/p_0_in [3]),
        .O(\r7/p_0_out [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[19]_i_1__6 
       (.I0(\r8/t0/t1/p_1_in [3]),
        .I1(\r8/t2/t3/p_0_in [3]),
        .I2(\r8/t1/t2/p_1_in [3]),
        .I3(\r8/t1/t2/p_0_in [3]),
        .I4(k7b[19]),
        .I5(\r8/t3/t0/p_0_in [3]),
        .O(\r8/p_0_out [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[19]_i_1__7 
       (.I0(\r9/t0/t1/p_1_in [3]),
        .I1(\r9/t2/t3/p_0_in [3]),
        .I2(\r9/t1/t2/p_1_in [3]),
        .I3(\r9/t1/t2/p_0_in [3]),
        .I4(k8b[19]),
        .I5(\r9/t3/t0/p_0_in [3]),
        .O(\r9/p_0_out [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair355" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[19]_i_1__8 
       (.I0(\a10/k3a [19]),
        .I1(\a10/k4a [19]),
        .I2(\rf/p_0_in [19]),
        .O(\rf/p_4_out [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[1]_i_1 
       (.I0(\r1/t0/t1/p_0_in [1]),
        .I1(\r1/t2/t3/p_1_in [1]),
        .I2(\r1/t1/t2/p_0_in [1]),
        .I3(k0b[1]),
        .I4(\r1/t3/t0/p_1_in [1]),
        .I5(\r1/t3/t0/p_0_in [1]),
        .O(\r1/p_0_out [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[1]_i_1__0 
       (.I0(\r2/t0/t1/p_0_in [1]),
        .I1(\r2/t2/t3/p_1_in [1]),
        .I2(\r2/t1/t2/p_0_in [1]),
        .I3(k1b[1]),
        .I4(\r2/t3/t0/p_1_in [1]),
        .I5(\r2/t3/t0/p_0_in [1]),
        .O(\r2/p_0_out [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[1]_i_1__1 
       (.I0(\r3/t0/t1/p_0_in [1]),
        .I1(\r3/t2/t3/p_1_in [1]),
        .I2(\r3/t1/t2/p_0_in [1]),
        .I3(k2b[1]),
        .I4(\r3/t3/t0/p_1_in [1]),
        .I5(\r3/t3/t0/p_0_in [1]),
        .O(\r3/p_0_out [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[1]_i_1__2 
       (.I0(\r4/t0/t1/p_0_in [1]),
        .I1(\r4/t2/t3/p_1_in [1]),
        .I2(\r4/t1/t2/p_0_in [1]),
        .I3(k3b[1]),
        .I4(\r4/t3/t0/p_1_in [1]),
        .I5(\r4/t3/t0/p_0_in [1]),
        .O(\r4/p_0_out [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[1]_i_1__3 
       (.I0(\r5/t0/t1/p_0_in [1]),
        .I1(\r5/t2/t3/p_1_in [1]),
        .I2(\r5/t1/t2/p_0_in [1]),
        .I3(k4b[1]),
        .I4(\r5/t3/t0/p_1_in [1]),
        .I5(\r5/t3/t0/p_0_in [1]),
        .O(\r5/p_0_out [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[1]_i_1__4 
       (.I0(\r6/t0/t1/p_0_in [1]),
        .I1(\r6/t2/t3/p_1_in [1]),
        .I2(\r6/t1/t2/p_0_in [1]),
        .I3(k5b[1]),
        .I4(\r6/t3/t0/p_1_in [1]),
        .I5(\r6/t3/t0/p_0_in [1]),
        .O(\r6/p_0_out [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[1]_i_1__5 
       (.I0(\r7/t0/t1/p_0_in [1]),
        .I1(\r7/t2/t3/p_1_in [1]),
        .I2(\r7/t1/t2/p_0_in [1]),
        .I3(k6b[1]),
        .I4(\r7/t3/t0/p_1_in [1]),
        .I5(\r7/t3/t0/p_0_in [1]),
        .O(\r7/p_0_out [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[1]_i_1__6 
       (.I0(\r8/t0/t1/p_0_in [1]),
        .I1(\r8/t2/t3/p_1_in [1]),
        .I2(\r8/t1/t2/p_0_in [1]),
        .I3(k7b[1]),
        .I4(\r8/t3/t0/p_1_in [1]),
        .I5(\r8/t3/t0/p_0_in [1]),
        .O(\r8/p_0_out [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[1]_i_1__7 
       (.I0(\r9/t0/t1/p_0_in [1]),
        .I1(\r9/t2/t3/p_1_in [1]),
        .I2(\r9/t1/t2/p_0_in [1]),
        .I3(k8b[1]),
        .I4(\r9/t3/t0/p_1_in [1]),
        .I5(\r9/t3/t0/p_0_in [1]),
        .O(\r9/p_0_out [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair341" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[1]_i_1__8 
       (.I0(\a10/k3a [1]),
        .I1(\a10/k4a [1]),
        .I2(\rf/p_0_in [1]),
        .O(\rf/p_4_out [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[20]_i_1 
       (.I0(\r1/t0/t1/p_1_in [4]),
        .I1(\r1/t2/t3/p_0_in [4]),
        .I2(\r1/t1/t2/p_1_in [4]),
        .I3(\r1/t1/t2/p_0_in [4]),
        .I4(k0b[20]),
        .I5(\r1/t3/t0/p_0_in [4]),
        .O(\r1/p_0_out [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[20]_i_1__0 
       (.I0(\r2/t0/t1/p_1_in [4]),
        .I1(\r2/t2/t3/p_0_in [4]),
        .I2(\r2/t1/t2/p_1_in [4]),
        .I3(\r2/t1/t2/p_0_in [4]),
        .I4(k1b[20]),
        .I5(\r2/t3/t0/p_0_in [4]),
        .O(\r2/p_0_out [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[20]_i_1__1 
       (.I0(\r3/t0/t1/p_1_in [4]),
        .I1(\r3/t2/t3/p_0_in [4]),
        .I2(\r3/t1/t2/p_1_in [4]),
        .I3(\r3/t1/t2/p_0_in [4]),
        .I4(k2b[20]),
        .I5(\r3/t3/t0/p_0_in [4]),
        .O(\r3/p_0_out [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[20]_i_1__2 
       (.I0(\r4/t0/t1/p_1_in [4]),
        .I1(\r4/t2/t3/p_0_in [4]),
        .I2(\r4/t1/t2/p_1_in [4]),
        .I3(\r4/t1/t2/p_0_in [4]),
        .I4(k3b[20]),
        .I5(\r4/t3/t0/p_0_in [4]),
        .O(\r4/p_0_out [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[20]_i_1__3 
       (.I0(\r5/t0/t1/p_1_in [4]),
        .I1(\r5/t2/t3/p_0_in [4]),
        .I2(\r5/t1/t2/p_1_in [4]),
        .I3(\r5/t1/t2/p_0_in [4]),
        .I4(k4b[20]),
        .I5(\r5/t3/t0/p_0_in [4]),
        .O(\r5/p_0_out [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[20]_i_1__4 
       (.I0(\r6/t0/t1/p_1_in [4]),
        .I1(\r6/t2/t3/p_0_in [4]),
        .I2(\r6/t1/t2/p_1_in [4]),
        .I3(\r6/t1/t2/p_0_in [4]),
        .I4(k5b[20]),
        .I5(\r6/t3/t0/p_0_in [4]),
        .O(\r6/p_0_out [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[20]_i_1__5 
       (.I0(\r7/t0/t1/p_1_in [4]),
        .I1(\r7/t2/t3/p_0_in [4]),
        .I2(\r7/t1/t2/p_1_in [4]),
        .I3(\r7/t1/t2/p_0_in [4]),
        .I4(k6b[20]),
        .I5(\r7/t3/t0/p_0_in [4]),
        .O(\r7/p_0_out [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[20]_i_1__6 
       (.I0(\r8/t0/t1/p_1_in [4]),
        .I1(\r8/t2/t3/p_0_in [4]),
        .I2(\r8/t1/t2/p_1_in [4]),
        .I3(\r8/t1/t2/p_0_in [4]),
        .I4(k7b[20]),
        .I5(\r8/t3/t0/p_0_in [4]),
        .O(\r8/p_0_out [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[20]_i_1__7 
       (.I0(\r9/t0/t1/p_1_in [4]),
        .I1(\r9/t2/t3/p_0_in [4]),
        .I2(\r9/t1/t2/p_1_in [4]),
        .I3(\r9/t1/t2/p_0_in [4]),
        .I4(k8b[20]),
        .I5(\r9/t3/t0/p_0_in [4]),
        .O(\r9/p_0_out [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair354" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[20]_i_1__8 
       (.I0(\a10/k3a [20]),
        .I1(\a10/k4a [20]),
        .I2(\rf/p_0_in [20]),
        .O(\rf/p_4_out [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[21]_i_1 
       (.I0(\r1/t0/t1/p_1_in [5]),
        .I1(\r1/t2/t3/p_0_in [5]),
        .I2(\r1/t1/t2/p_1_in [5]),
        .I3(\r1/t1/t2/p_0_in [5]),
        .I4(k0b[21]),
        .I5(\r1/t3/t0/p_0_in [5]),
        .O(\r1/p_0_out [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[21]_i_1__0 
       (.I0(\r2/t0/t1/p_1_in [5]),
        .I1(\r2/t2/t3/p_0_in [5]),
        .I2(\r2/t1/t2/p_1_in [5]),
        .I3(\r2/t1/t2/p_0_in [5]),
        .I4(k1b[21]),
        .I5(\r2/t3/t0/p_0_in [5]),
        .O(\r2/p_0_out [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[21]_i_1__1 
       (.I0(\r3/t0/t1/p_1_in [5]),
        .I1(\r3/t2/t3/p_0_in [5]),
        .I2(\r3/t1/t2/p_1_in [5]),
        .I3(\r3/t1/t2/p_0_in [5]),
        .I4(k2b[21]),
        .I5(\r3/t3/t0/p_0_in [5]),
        .O(\r3/p_0_out [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[21]_i_1__2 
       (.I0(\r4/t0/t1/p_1_in [5]),
        .I1(\r4/t2/t3/p_0_in [5]),
        .I2(\r4/t1/t2/p_1_in [5]),
        .I3(\r4/t1/t2/p_0_in [5]),
        .I4(k3b[21]),
        .I5(\r4/t3/t0/p_0_in [5]),
        .O(\r4/p_0_out [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[21]_i_1__3 
       (.I0(\r5/t0/t1/p_1_in [5]),
        .I1(\r5/t2/t3/p_0_in [5]),
        .I2(\r5/t1/t2/p_1_in [5]),
        .I3(\r5/t1/t2/p_0_in [5]),
        .I4(k4b[21]),
        .I5(\r5/t3/t0/p_0_in [5]),
        .O(\r5/p_0_out [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[21]_i_1__4 
       (.I0(\r6/t0/t1/p_1_in [5]),
        .I1(\r6/t2/t3/p_0_in [5]),
        .I2(\r6/t1/t2/p_1_in [5]),
        .I3(\r6/t1/t2/p_0_in [5]),
        .I4(k5b[21]),
        .I5(\r6/t3/t0/p_0_in [5]),
        .O(\r6/p_0_out [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[21]_i_1__5 
       (.I0(\r7/t0/t1/p_1_in [5]),
        .I1(\r7/t2/t3/p_0_in [5]),
        .I2(\r7/t1/t2/p_1_in [5]),
        .I3(\r7/t1/t2/p_0_in [5]),
        .I4(k6b[21]),
        .I5(\r7/t3/t0/p_0_in [5]),
        .O(\r7/p_0_out [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[21]_i_1__6 
       (.I0(\r8/t0/t1/p_1_in [5]),
        .I1(\r8/t2/t3/p_0_in [5]),
        .I2(\r8/t1/t2/p_1_in [5]),
        .I3(\r8/t1/t2/p_0_in [5]),
        .I4(k7b[21]),
        .I5(\r8/t3/t0/p_0_in [5]),
        .O(\r8/p_0_out [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[21]_i_1__7 
       (.I0(\r9/t0/t1/p_1_in [5]),
        .I1(\r9/t2/t3/p_0_in [5]),
        .I2(\r9/t1/t2/p_1_in [5]),
        .I3(\r9/t1/t2/p_0_in [5]),
        .I4(k8b[21]),
        .I5(\r9/t3/t0/p_0_in [5]),
        .O(\r9/p_0_out [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair353" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[21]_i_1__8 
       (.I0(\a10/k3a [21]),
        .I1(\a10/k4a [21]),
        .I2(\rf/p_0_in [21]),
        .O(\rf/p_4_out [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[22]_i_1 
       (.I0(\r1/t0/t1/p_1_in [6]),
        .I1(\r1/t2/t3/p_0_in [6]),
        .I2(\r1/t1/t2/p_1_in [6]),
        .I3(\r1/t1/t2/p_0_in [6]),
        .I4(k0b[22]),
        .I5(\r1/t3/t0/p_0_in [6]),
        .O(\r1/p_0_out [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[22]_i_1__0 
       (.I0(\r2/t0/t1/p_1_in [6]),
        .I1(\r2/t2/t3/p_0_in [6]),
        .I2(\r2/t1/t2/p_1_in [6]),
        .I3(\r2/t1/t2/p_0_in [6]),
        .I4(k1b[22]),
        .I5(\r2/t3/t0/p_0_in [6]),
        .O(\r2/p_0_out [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[22]_i_1__1 
       (.I0(\r3/t0/t1/p_1_in [6]),
        .I1(\r3/t2/t3/p_0_in [6]),
        .I2(\r3/t1/t2/p_1_in [6]),
        .I3(\r3/t1/t2/p_0_in [6]),
        .I4(k2b[22]),
        .I5(\r3/t3/t0/p_0_in [6]),
        .O(\r3/p_0_out [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[22]_i_1__2 
       (.I0(\r4/t0/t1/p_1_in [6]),
        .I1(\r4/t2/t3/p_0_in [6]),
        .I2(\r4/t1/t2/p_1_in [6]),
        .I3(\r4/t1/t2/p_0_in [6]),
        .I4(k3b[22]),
        .I5(\r4/t3/t0/p_0_in [6]),
        .O(\r4/p_0_out [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[22]_i_1__3 
       (.I0(\r5/t0/t1/p_1_in [6]),
        .I1(\r5/t2/t3/p_0_in [6]),
        .I2(\r5/t1/t2/p_1_in [6]),
        .I3(\r5/t1/t2/p_0_in [6]),
        .I4(k4b[22]),
        .I5(\r5/t3/t0/p_0_in [6]),
        .O(\r5/p_0_out [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[22]_i_1__4 
       (.I0(\r6/t0/t1/p_1_in [6]),
        .I1(\r6/t2/t3/p_0_in [6]),
        .I2(\r6/t1/t2/p_1_in [6]),
        .I3(\r6/t1/t2/p_0_in [6]),
        .I4(k5b[22]),
        .I5(\r6/t3/t0/p_0_in [6]),
        .O(\r6/p_0_out [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[22]_i_1__5 
       (.I0(\r7/t0/t1/p_1_in [6]),
        .I1(\r7/t2/t3/p_0_in [6]),
        .I2(\r7/t1/t2/p_1_in [6]),
        .I3(\r7/t1/t2/p_0_in [6]),
        .I4(k6b[22]),
        .I5(\r7/t3/t0/p_0_in [6]),
        .O(\r7/p_0_out [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[22]_i_1__6 
       (.I0(\r8/t0/t1/p_1_in [6]),
        .I1(\r8/t2/t3/p_0_in [6]),
        .I2(\r8/t1/t2/p_1_in [6]),
        .I3(\r8/t1/t2/p_0_in [6]),
        .I4(k7b[22]),
        .I5(\r8/t3/t0/p_0_in [6]),
        .O(\r8/p_0_out [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[22]_i_1__7 
       (.I0(\r9/t0/t1/p_1_in [6]),
        .I1(\r9/t2/t3/p_0_in [6]),
        .I2(\r9/t1/t2/p_1_in [6]),
        .I3(\r9/t1/t2/p_0_in [6]),
        .I4(k8b[22]),
        .I5(\r9/t3/t0/p_0_in [6]),
        .O(\r9/p_0_out [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair352" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[22]_i_1__8 
       (.I0(\a10/k3a [22]),
        .I1(\a10/k4a [22]),
        .I2(\rf/p_0_in [22]),
        .O(\rf/p_4_out [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[23]_i_1 
       (.I0(\r1/t0/t1/p_1_in [7]),
        .I1(\r1/t2/t3/p_0_in [7]),
        .I2(\r1/t1/t2/p_1_in [7]),
        .I3(\r1/t1/t2/p_0_in [7]),
        .I4(k0b[23]),
        .I5(\r1/t3/t0/p_0_in [7]),
        .O(\r1/p_0_out [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[23]_i_1__0 
       (.I0(\r2/t0/t1/p_1_in [7]),
        .I1(\r2/t2/t3/p_0_in [7]),
        .I2(\r2/t1/t2/p_1_in [7]),
        .I3(\r2/t1/t2/p_0_in [7]),
        .I4(k1b[23]),
        .I5(\r2/t3/t0/p_0_in [7]),
        .O(\r2/p_0_out [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[23]_i_1__1 
       (.I0(\r3/t0/t1/p_1_in [7]),
        .I1(\r3/t2/t3/p_0_in [7]),
        .I2(\r3/t1/t2/p_1_in [7]),
        .I3(\r3/t1/t2/p_0_in [7]),
        .I4(k2b[23]),
        .I5(\r3/t3/t0/p_0_in [7]),
        .O(\r3/p_0_out [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[23]_i_1__2 
       (.I0(\r4/t0/t1/p_1_in [7]),
        .I1(\r4/t2/t3/p_0_in [7]),
        .I2(\r4/t1/t2/p_1_in [7]),
        .I3(\r4/t1/t2/p_0_in [7]),
        .I4(k3b[23]),
        .I5(\r4/t3/t0/p_0_in [7]),
        .O(\r4/p_0_out [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[23]_i_1__3 
       (.I0(\r5/t0/t1/p_1_in [7]),
        .I1(\r5/t2/t3/p_0_in [7]),
        .I2(\r5/t1/t2/p_1_in [7]),
        .I3(\r5/t1/t2/p_0_in [7]),
        .I4(k4b[23]),
        .I5(\r5/t3/t0/p_0_in [7]),
        .O(\r5/p_0_out [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[23]_i_1__4 
       (.I0(\r6/t0/t1/p_1_in [7]),
        .I1(\r6/t2/t3/p_0_in [7]),
        .I2(\r6/t1/t2/p_1_in [7]),
        .I3(\r6/t1/t2/p_0_in [7]),
        .I4(k5b[23]),
        .I5(\r6/t3/t0/p_0_in [7]),
        .O(\r6/p_0_out [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[23]_i_1__5 
       (.I0(\r7/t0/t1/p_1_in [7]),
        .I1(\r7/t2/t3/p_0_in [7]),
        .I2(\r7/t1/t2/p_1_in [7]),
        .I3(\r7/t1/t2/p_0_in [7]),
        .I4(k6b[23]),
        .I5(\r7/t3/t0/p_0_in [7]),
        .O(\r7/p_0_out [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[23]_i_1__6 
       (.I0(\r8/t0/t1/p_1_in [7]),
        .I1(\r8/t2/t3/p_0_in [7]),
        .I2(\r8/t1/t2/p_1_in [7]),
        .I3(\r8/t1/t2/p_0_in [7]),
        .I4(k7b[23]),
        .I5(\r8/t3/t0/p_0_in [7]),
        .O(\r8/p_0_out [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[23]_i_1__7 
       (.I0(\r9/t0/t1/p_1_in [7]),
        .I1(\r9/t2/t3/p_0_in [7]),
        .I2(\r9/t1/t2/p_1_in [7]),
        .I3(\r9/t1/t2/p_0_in [7]),
        .I4(k8b[23]),
        .I5(\r9/t3/t0/p_0_in [7]),
        .O(\r9/p_0_out [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair351" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[23]_i_1__8 
       (.I0(\a10/k3a [23]),
        .I1(\a10/k4a [23]),
        .I2(\rf/p_0_in [23]),
        .O(\rf/p_4_out [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[24]_i_1 
       (.I0(\r1/t0/t1/p_1_in [0]),
        .I1(\r1/t0/t1/p_0_in [0]),
        .I2(\r1/t2/t3/p_0_in [0]),
        .I3(\r1/t1/t2/p_0_in [0]),
        .I4(k0b[24]),
        .I5(\r1/t3/t0/p_1_in [0]),
        .O(\r1/p_0_out [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[24]_i_1__0 
       (.I0(\r2/t0/t1/p_1_in [0]),
        .I1(\r2/t0/t1/p_0_in [0]),
        .I2(\r2/t2/t3/p_0_in [0]),
        .I3(\r2/t1/t2/p_0_in [0]),
        .I4(k1b[24]),
        .I5(\r2/t3/t0/p_1_in [0]),
        .O(\r2/p_0_out [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[24]_i_1__1 
       (.I0(\r3/t0/t1/p_1_in [0]),
        .I1(\r3/t0/t1/p_0_in [0]),
        .I2(\r3/t2/t3/p_0_in [0]),
        .I3(\r3/t1/t2/p_0_in [0]),
        .I4(k2b[24]),
        .I5(\r3/t3/t0/p_1_in [0]),
        .O(\r3/p_0_out [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[24]_i_1__2 
       (.I0(\r4/t0/t1/p_1_in [0]),
        .I1(\r4/t0/t1/p_0_in [0]),
        .I2(\r4/t2/t3/p_0_in [0]),
        .I3(\r4/t1/t2/p_0_in [0]),
        .I4(k3b[24]),
        .I5(\r4/t3/t0/p_1_in [0]),
        .O(\r4/p_0_out [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[24]_i_1__3 
       (.I0(\r5/t0/t1/p_1_in [0]),
        .I1(\r5/t0/t1/p_0_in [0]),
        .I2(\r5/t2/t3/p_0_in [0]),
        .I3(\r5/t1/t2/p_0_in [0]),
        .I4(k4b[24]),
        .I5(\r5/t3/t0/p_1_in [0]),
        .O(\r5/p_0_out [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[24]_i_1__4 
       (.I0(\r6/t0/t1/p_1_in [0]),
        .I1(\r6/t0/t1/p_0_in [0]),
        .I2(\r6/t2/t3/p_0_in [0]),
        .I3(\r6/t1/t2/p_0_in [0]),
        .I4(k5b[24]),
        .I5(\r6/t3/t0/p_1_in [0]),
        .O(\r6/p_0_out [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[24]_i_1__5 
       (.I0(\r7/t0/t1/p_1_in [0]),
        .I1(\r7/t0/t1/p_0_in [0]),
        .I2(\r7/t2/t3/p_0_in [0]),
        .I3(\r7/t1/t2/p_0_in [0]),
        .I4(k6b[24]),
        .I5(\r7/t3/t0/p_1_in [0]),
        .O(\r7/p_0_out [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[24]_i_1__6 
       (.I0(\r8/t0/t1/p_1_in [0]),
        .I1(\r8/t0/t1/p_0_in [0]),
        .I2(\r8/t2/t3/p_0_in [0]),
        .I3(\r8/t1/t2/p_0_in [0]),
        .I4(k7b[24]),
        .I5(\r8/t3/t0/p_1_in [0]),
        .O(\r8/p_0_out [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[24]_i_1__7 
       (.I0(\r9/t0/t1/p_1_in [0]),
        .I1(\r9/t0/t1/p_0_in [0]),
        .I2(\r9/t2/t3/p_0_in [0]),
        .I3(\r9/t1/t2/p_0_in [0]),
        .I4(k8b[24]),
        .I5(\r9/t3/t0/p_1_in [0]),
        .O(\r9/p_0_out [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair325" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[24]_i_1__8 
       (.I0(\a10/k3a [24]),
        .I1(\a10/k4a [24]),
        .I2(\rf/p_0_in [24]),
        .O(\rf/p_4_out [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[25]_i_1 
       (.I0(\r1/t0/t1/p_1_in [1]),
        .I1(\r1/t0/t1/p_0_in [1]),
        .I2(\r1/t2/t3/p_0_in [1]),
        .I3(\r1/t1/t2/p_0_in [1]),
        .I4(k0b[25]),
        .I5(\r1/t3/t0/p_1_in [1]),
        .O(\r1/p_0_out [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[25]_i_1__0 
       (.I0(\r2/t0/t1/p_1_in [1]),
        .I1(\r2/t0/t1/p_0_in [1]),
        .I2(\r2/t2/t3/p_0_in [1]),
        .I3(\r2/t1/t2/p_0_in [1]),
        .I4(k1b[25]),
        .I5(\r2/t3/t0/p_1_in [1]),
        .O(\r2/p_0_out [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[25]_i_1__1 
       (.I0(\r3/t0/t1/p_1_in [1]),
        .I1(\r3/t0/t1/p_0_in [1]),
        .I2(\r3/t2/t3/p_0_in [1]),
        .I3(\r3/t1/t2/p_0_in [1]),
        .I4(k2b[25]),
        .I5(\r3/t3/t0/p_1_in [1]),
        .O(\r3/p_0_out [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[25]_i_1__2 
       (.I0(\r4/t0/t1/p_1_in [1]),
        .I1(\r4/t0/t1/p_0_in [1]),
        .I2(\r4/t2/t3/p_0_in [1]),
        .I3(\r4/t1/t2/p_0_in [1]),
        .I4(k3b[25]),
        .I5(\r4/t3/t0/p_1_in [1]),
        .O(\r4/p_0_out [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[25]_i_1__3 
       (.I0(\r5/t0/t1/p_1_in [1]),
        .I1(\r5/t0/t1/p_0_in [1]),
        .I2(\r5/t2/t3/p_0_in [1]),
        .I3(\r5/t1/t2/p_0_in [1]),
        .I4(k4b[25]),
        .I5(\r5/t3/t0/p_1_in [1]),
        .O(\r5/p_0_out [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[25]_i_1__4 
       (.I0(\r6/t0/t1/p_1_in [1]),
        .I1(\r6/t0/t1/p_0_in [1]),
        .I2(\r6/t2/t3/p_0_in [1]),
        .I3(\r6/t1/t2/p_0_in [1]),
        .I4(k5b[25]),
        .I5(\r6/t3/t0/p_1_in [1]),
        .O(\r6/p_0_out [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[25]_i_1__5 
       (.I0(\r7/t0/t1/p_1_in [1]),
        .I1(\r7/t0/t1/p_0_in [1]),
        .I2(\r7/t2/t3/p_0_in [1]),
        .I3(\r7/t1/t2/p_0_in [1]),
        .I4(k6b[25]),
        .I5(\r7/t3/t0/p_1_in [1]),
        .O(\r7/p_0_out [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[25]_i_1__6 
       (.I0(\r8/t0/t1/p_1_in [1]),
        .I1(\r8/t0/t1/p_0_in [1]),
        .I2(\r8/t2/t3/p_0_in [1]),
        .I3(\r8/t1/t2/p_0_in [1]),
        .I4(k7b[25]),
        .I5(\r8/t3/t0/p_1_in [1]),
        .O(\r8/p_0_out [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[25]_i_1__7 
       (.I0(\r9/t0/t1/p_1_in [1]),
        .I1(\r9/t0/t1/p_0_in [1]),
        .I2(\r9/t2/t3/p_0_in [1]),
        .I3(\r9/t1/t2/p_0_in [1]),
        .I4(k8b[25]),
        .I5(\r9/t3/t0/p_1_in [1]),
        .O(\r9/p_0_out [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair322" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[25]_i_1__8 
       (.I0(\a10/k3a [25]),
        .I1(\a10/k4a [25]),
        .I2(\rf/p_0_in [25]),
        .O(\rf/p_4_out [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[26]_i_1 
       (.I0(\r1/t0/t1/p_1_in [2]),
        .I1(\r1/t0/t1/p_0_in [2]),
        .I2(\r1/t2/t3/p_0_in [2]),
        .I3(\r1/t1/t2/p_0_in [2]),
        .I4(k0b[26]),
        .I5(\r1/t3/t0/p_1_in [2]),
        .O(\r1/p_0_out [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[26]_i_1__0 
       (.I0(\r2/t0/t1/p_1_in [2]),
        .I1(\r2/t0/t1/p_0_in [2]),
        .I2(\r2/t2/t3/p_0_in [2]),
        .I3(\r2/t1/t2/p_0_in [2]),
        .I4(k1b[26]),
        .I5(\r2/t3/t0/p_1_in [2]),
        .O(\r2/p_0_out [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[26]_i_1__1 
       (.I0(\r3/t0/t1/p_1_in [2]),
        .I1(\r3/t0/t1/p_0_in [2]),
        .I2(\r3/t2/t3/p_0_in [2]),
        .I3(\r3/t1/t2/p_0_in [2]),
        .I4(k2b[26]),
        .I5(\r3/t3/t0/p_1_in [2]),
        .O(\r3/p_0_out [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[26]_i_1__2 
       (.I0(\r4/t0/t1/p_1_in [2]),
        .I1(\r4/t0/t1/p_0_in [2]),
        .I2(\r4/t2/t3/p_0_in [2]),
        .I3(\r4/t1/t2/p_0_in [2]),
        .I4(k3b[26]),
        .I5(\r4/t3/t0/p_1_in [2]),
        .O(\r4/p_0_out [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[26]_i_1__3 
       (.I0(\r5/t0/t1/p_1_in [2]),
        .I1(\r5/t0/t1/p_0_in [2]),
        .I2(\r5/t2/t3/p_0_in [2]),
        .I3(\r5/t1/t2/p_0_in [2]),
        .I4(k4b[26]),
        .I5(\r5/t3/t0/p_1_in [2]),
        .O(\r5/p_0_out [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[26]_i_1__4 
       (.I0(\r6/t0/t1/p_1_in [2]),
        .I1(\r6/t0/t1/p_0_in [2]),
        .I2(\r6/t2/t3/p_0_in [2]),
        .I3(\r6/t1/t2/p_0_in [2]),
        .I4(k5b[26]),
        .I5(\r6/t3/t0/p_1_in [2]),
        .O(\r6/p_0_out [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[26]_i_1__5 
       (.I0(\r7/t0/t1/p_1_in [2]),
        .I1(\r7/t0/t1/p_0_in [2]),
        .I2(\r7/t2/t3/p_0_in [2]),
        .I3(\r7/t1/t2/p_0_in [2]),
        .I4(k6b[26]),
        .I5(\r7/t3/t0/p_1_in [2]),
        .O(\r7/p_0_out [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[26]_i_1__6 
       (.I0(\r8/t0/t1/p_1_in [2]),
        .I1(\r8/t0/t1/p_0_in [2]),
        .I2(\r8/t2/t3/p_0_in [2]),
        .I3(\r8/t1/t2/p_0_in [2]),
        .I4(k7b[26]),
        .I5(\r8/t3/t0/p_1_in [2]),
        .O(\r8/p_0_out [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[26]_i_1__7 
       (.I0(\r9/t0/t1/p_1_in [2]),
        .I1(\r9/t0/t1/p_0_in [2]),
        .I2(\r9/t2/t3/p_0_in [2]),
        .I3(\r9/t1/t2/p_0_in [2]),
        .I4(k8b[26]),
        .I5(\r9/t3/t0/p_1_in [2]),
        .O(\r9/p_0_out [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair327" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[26]_i_1__8 
       (.I0(\a10/k3a [26]),
        .I1(\a10/k4a [26]),
        .I2(\rf/p_0_in [26]),
        .O(\rf/p_4_out [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[27]_i_1 
       (.I0(\r1/t0/t1/p_1_in [3]),
        .I1(\r1/t0/t1/p_0_in [3]),
        .I2(\r1/t2/t3/p_0_in [3]),
        .I3(\r1/t1/t2/p_0_in [3]),
        .I4(k0b[27]),
        .I5(\r1/t3/t0/p_1_in [3]),
        .O(\r1/p_0_out [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[27]_i_1__0 
       (.I0(\r2/t0/t1/p_1_in [3]),
        .I1(\r2/t0/t1/p_0_in [3]),
        .I2(\r2/t2/t3/p_0_in [3]),
        .I3(\r2/t1/t2/p_0_in [3]),
        .I4(k1b[27]),
        .I5(\r2/t3/t0/p_1_in [3]),
        .O(\r2/p_0_out [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[27]_i_1__1 
       (.I0(\r3/t0/t1/p_1_in [3]),
        .I1(\r3/t0/t1/p_0_in [3]),
        .I2(\r3/t2/t3/p_0_in [3]),
        .I3(\r3/t1/t2/p_0_in [3]),
        .I4(k2b[27]),
        .I5(\r3/t3/t0/p_1_in [3]),
        .O(\r3/p_0_out [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[27]_i_1__2 
       (.I0(\r4/t0/t1/p_1_in [3]),
        .I1(\r4/t0/t1/p_0_in [3]),
        .I2(\r4/t2/t3/p_0_in [3]),
        .I3(\r4/t1/t2/p_0_in [3]),
        .I4(k3b[27]),
        .I5(\r4/t3/t0/p_1_in [3]),
        .O(\r4/p_0_out [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[27]_i_1__3 
       (.I0(\r5/t0/t1/p_1_in [3]),
        .I1(\r5/t0/t1/p_0_in [3]),
        .I2(\r5/t2/t3/p_0_in [3]),
        .I3(\r5/t1/t2/p_0_in [3]),
        .I4(k4b[27]),
        .I5(\r5/t3/t0/p_1_in [3]),
        .O(\r5/p_0_out [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[27]_i_1__4 
       (.I0(\r6/t0/t1/p_1_in [3]),
        .I1(\r6/t0/t1/p_0_in [3]),
        .I2(\r6/t2/t3/p_0_in [3]),
        .I3(\r6/t1/t2/p_0_in [3]),
        .I4(k5b[27]),
        .I5(\r6/t3/t0/p_1_in [3]),
        .O(\r6/p_0_out [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[27]_i_1__5 
       (.I0(\r7/t0/t1/p_1_in [3]),
        .I1(\r7/t0/t1/p_0_in [3]),
        .I2(\r7/t2/t3/p_0_in [3]),
        .I3(\r7/t1/t2/p_0_in [3]),
        .I4(k6b[27]),
        .I5(\r7/t3/t0/p_1_in [3]),
        .O(\r7/p_0_out [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[27]_i_1__6 
       (.I0(\r8/t0/t1/p_1_in [3]),
        .I1(\r8/t0/t1/p_0_in [3]),
        .I2(\r8/t2/t3/p_0_in [3]),
        .I3(\r8/t1/t2/p_0_in [3]),
        .I4(k7b[27]),
        .I5(\r8/t3/t0/p_1_in [3]),
        .O(\r8/p_0_out [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[27]_i_1__7 
       (.I0(\r9/t0/t1/p_1_in [3]),
        .I1(\r9/t0/t1/p_0_in [3]),
        .I2(\r9/t2/t3/p_0_in [3]),
        .I3(\r9/t1/t2/p_0_in [3]),
        .I4(k8b[27]),
        .I5(\r9/t3/t0/p_1_in [3]),
        .O(\r9/p_0_out [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair326" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[27]_i_1__8 
       (.I0(\a10/k3a [27]),
        .I1(\a10/k4a [27]),
        .I2(\rf/p_0_in [27]),
        .O(\rf/p_4_out [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[28]_i_1 
       (.I0(\r1/t0/t1/p_1_in [4]),
        .I1(\r1/t0/t1/p_0_in [4]),
        .I2(\r1/t2/t3/p_0_in [4]),
        .I3(\r1/t1/t2/p_0_in [4]),
        .I4(k0b[28]),
        .I5(\r1/t3/t0/p_1_in [4]),
        .O(\r1/p_0_out [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[28]_i_1__0 
       (.I0(\r2/t0/t1/p_1_in [4]),
        .I1(\r2/t0/t1/p_0_in [4]),
        .I2(\r2/t2/t3/p_0_in [4]),
        .I3(\r2/t1/t2/p_0_in [4]),
        .I4(k1b[28]),
        .I5(\r2/t3/t0/p_1_in [4]),
        .O(\r2/p_0_out [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[28]_i_1__1 
       (.I0(\r3/t0/t1/p_1_in [4]),
        .I1(\r3/t0/t1/p_0_in [4]),
        .I2(\r3/t2/t3/p_0_in [4]),
        .I3(\r3/t1/t2/p_0_in [4]),
        .I4(k2b[28]),
        .I5(\r3/t3/t0/p_1_in [4]),
        .O(\r3/p_0_out [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[28]_i_1__2 
       (.I0(\r4/t0/t1/p_1_in [4]),
        .I1(\r4/t0/t1/p_0_in [4]),
        .I2(\r4/t2/t3/p_0_in [4]),
        .I3(\r4/t1/t2/p_0_in [4]),
        .I4(k3b[28]),
        .I5(\r4/t3/t0/p_1_in [4]),
        .O(\r4/p_0_out [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[28]_i_1__3 
       (.I0(\r5/t0/t1/p_1_in [4]),
        .I1(\r5/t0/t1/p_0_in [4]),
        .I2(\r5/t2/t3/p_0_in [4]),
        .I3(\r5/t1/t2/p_0_in [4]),
        .I4(k4b[28]),
        .I5(\r5/t3/t0/p_1_in [4]),
        .O(\r5/p_0_out [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[28]_i_1__4 
       (.I0(\r6/t0/t1/p_1_in [4]),
        .I1(\r6/t0/t1/p_0_in [4]),
        .I2(\r6/t2/t3/p_0_in [4]),
        .I3(\r6/t1/t2/p_0_in [4]),
        .I4(k5b[28]),
        .I5(\r6/t3/t0/p_1_in [4]),
        .O(\r6/p_0_out [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[28]_i_1__5 
       (.I0(\r7/t0/t1/p_1_in [4]),
        .I1(\r7/t0/t1/p_0_in [4]),
        .I2(\r7/t2/t3/p_0_in [4]),
        .I3(\r7/t1/t2/p_0_in [4]),
        .I4(k6b[28]),
        .I5(\r7/t3/t0/p_1_in [4]),
        .O(\r7/p_0_out [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[28]_i_1__6 
       (.I0(\r8/t0/t1/p_1_in [4]),
        .I1(\r8/t0/t1/p_0_in [4]),
        .I2(\r8/t2/t3/p_0_in [4]),
        .I3(\r8/t1/t2/p_0_in [4]),
        .I4(k7b[28]),
        .I5(\r8/t3/t0/p_1_in [4]),
        .O(\r8/p_0_out [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[28]_i_1__7 
       (.I0(\r9/t0/t1/p_1_in [4]),
        .I1(\r9/t0/t1/p_0_in [4]),
        .I2(\r9/t2/t3/p_0_in [4]),
        .I3(\r9/t1/t2/p_0_in [4]),
        .I4(k8b[28]),
        .I5(\r9/t3/t0/p_1_in [4]),
        .O(\r9/p_0_out [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair320" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[28]_i_1__8 
       (.I0(\a10/k3a [28]),
        .I1(\a10/k4a [28]),
        .I2(\rf/p_0_in [28]),
        .O(\rf/p_4_out [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[29]_i_1 
       (.I0(\r1/t0/t1/p_1_in [5]),
        .I1(\r1/t0/t1/p_0_in [5]),
        .I2(\r1/t2/t3/p_0_in [5]),
        .I3(\r1/t1/t2/p_0_in [5]),
        .I4(k0b[29]),
        .I5(\r1/t3/t0/p_1_in [5]),
        .O(\r1/p_0_out [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[29]_i_1__0 
       (.I0(\r2/t0/t1/p_1_in [5]),
        .I1(\r2/t0/t1/p_0_in [5]),
        .I2(\r2/t2/t3/p_0_in [5]),
        .I3(\r2/t1/t2/p_0_in [5]),
        .I4(k1b[29]),
        .I5(\r2/t3/t0/p_1_in [5]),
        .O(\r2/p_0_out [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[29]_i_1__1 
       (.I0(\r3/t0/t1/p_1_in [5]),
        .I1(\r3/t0/t1/p_0_in [5]),
        .I2(\r3/t2/t3/p_0_in [5]),
        .I3(\r3/t1/t2/p_0_in [5]),
        .I4(k2b[29]),
        .I5(\r3/t3/t0/p_1_in [5]),
        .O(\r3/p_0_out [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[29]_i_1__2 
       (.I0(\r4/t0/t1/p_1_in [5]),
        .I1(\r4/t0/t1/p_0_in [5]),
        .I2(\r4/t2/t3/p_0_in [5]),
        .I3(\r4/t1/t2/p_0_in [5]),
        .I4(k3b[29]),
        .I5(\r4/t3/t0/p_1_in [5]),
        .O(\r4/p_0_out [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[29]_i_1__3 
       (.I0(\r5/t0/t1/p_1_in [5]),
        .I1(\r5/t0/t1/p_0_in [5]),
        .I2(\r5/t2/t3/p_0_in [5]),
        .I3(\r5/t1/t2/p_0_in [5]),
        .I4(k4b[29]),
        .I5(\r5/t3/t0/p_1_in [5]),
        .O(\r5/p_0_out [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[29]_i_1__4 
       (.I0(\r6/t0/t1/p_1_in [5]),
        .I1(\r6/t0/t1/p_0_in [5]),
        .I2(\r6/t2/t3/p_0_in [5]),
        .I3(\r6/t1/t2/p_0_in [5]),
        .I4(k5b[29]),
        .I5(\r6/t3/t0/p_1_in [5]),
        .O(\r6/p_0_out [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[29]_i_1__5 
       (.I0(\r7/t0/t1/p_1_in [5]),
        .I1(\r7/t0/t1/p_0_in [5]),
        .I2(\r7/t2/t3/p_0_in [5]),
        .I3(\r7/t1/t2/p_0_in [5]),
        .I4(k6b[29]),
        .I5(\r7/t3/t0/p_1_in [5]),
        .O(\r7/p_0_out [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[29]_i_1__6 
       (.I0(\r8/t0/t1/p_1_in [5]),
        .I1(\r8/t0/t1/p_0_in [5]),
        .I2(\r8/t2/t3/p_0_in [5]),
        .I3(\r8/t1/t2/p_0_in [5]),
        .I4(k7b[29]),
        .I5(\r8/t3/t0/p_1_in [5]),
        .O(\r8/p_0_out [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[29]_i_1__7 
       (.I0(\r9/t0/t1/p_1_in [5]),
        .I1(\r9/t0/t1/p_0_in [5]),
        .I2(\r9/t2/t3/p_0_in [5]),
        .I3(\r9/t1/t2/p_0_in [5]),
        .I4(k8b[29]),
        .I5(\r9/t3/t0/p_1_in [5]),
        .O(\r9/p_0_out [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair321" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[29]_i_1__8 
       (.I0(\a10/k3a [29]),
        .I1(\a10/k4a [29]),
        .I2(\rf/p_0_in [29]),
        .O(\rf/p_4_out [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[2]_i_1 
       (.I0(\r1/t0/t1/p_0_in [2]),
        .I1(\r1/t2/t3/p_1_in [2]),
        .I2(\r1/t1/t2/p_0_in [2]),
        .I3(k0b[2]),
        .I4(\r1/t3/t0/p_1_in [2]),
        .I5(\r1/t3/t0/p_0_in [2]),
        .O(\r1/p_0_out [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[2]_i_1__0 
       (.I0(\r2/t0/t1/p_0_in [2]),
        .I1(\r2/t2/t3/p_1_in [2]),
        .I2(\r2/t1/t2/p_0_in [2]),
        .I3(k1b[2]),
        .I4(\r2/t3/t0/p_1_in [2]),
        .I5(\r2/t3/t0/p_0_in [2]),
        .O(\r2/p_0_out [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[2]_i_1__1 
       (.I0(\r3/t0/t1/p_0_in [2]),
        .I1(\r3/t2/t3/p_1_in [2]),
        .I2(\r3/t1/t2/p_0_in [2]),
        .I3(k2b[2]),
        .I4(\r3/t3/t0/p_1_in [2]),
        .I5(\r3/t3/t0/p_0_in [2]),
        .O(\r3/p_0_out [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[2]_i_1__2 
       (.I0(\r4/t0/t1/p_0_in [2]),
        .I1(\r4/t2/t3/p_1_in [2]),
        .I2(\r4/t1/t2/p_0_in [2]),
        .I3(k3b[2]),
        .I4(\r4/t3/t0/p_1_in [2]),
        .I5(\r4/t3/t0/p_0_in [2]),
        .O(\r4/p_0_out [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[2]_i_1__3 
       (.I0(\r5/t0/t1/p_0_in [2]),
        .I1(\r5/t2/t3/p_1_in [2]),
        .I2(\r5/t1/t2/p_0_in [2]),
        .I3(k4b[2]),
        .I4(\r5/t3/t0/p_1_in [2]),
        .I5(\r5/t3/t0/p_0_in [2]),
        .O(\r5/p_0_out [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[2]_i_1__4 
       (.I0(\r6/t0/t1/p_0_in [2]),
        .I1(\r6/t2/t3/p_1_in [2]),
        .I2(\r6/t1/t2/p_0_in [2]),
        .I3(k5b[2]),
        .I4(\r6/t3/t0/p_1_in [2]),
        .I5(\r6/t3/t0/p_0_in [2]),
        .O(\r6/p_0_out [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[2]_i_1__5 
       (.I0(\r7/t0/t1/p_0_in [2]),
        .I1(\r7/t2/t3/p_1_in [2]),
        .I2(\r7/t1/t2/p_0_in [2]),
        .I3(k6b[2]),
        .I4(\r7/t3/t0/p_1_in [2]),
        .I5(\r7/t3/t0/p_0_in [2]),
        .O(\r7/p_0_out [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[2]_i_1__6 
       (.I0(\r8/t0/t1/p_0_in [2]),
        .I1(\r8/t2/t3/p_1_in [2]),
        .I2(\r8/t1/t2/p_0_in [2]),
        .I3(k7b[2]),
        .I4(\r8/t3/t0/p_1_in [2]),
        .I5(\r8/t3/t0/p_0_in [2]),
        .O(\r8/p_0_out [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[2]_i_1__7 
       (.I0(\r9/t0/t1/p_0_in [2]),
        .I1(\r9/t2/t3/p_1_in [2]),
        .I2(\r9/t1/t2/p_0_in [2]),
        .I3(k8b[2]),
        .I4(\r9/t3/t0/p_1_in [2]),
        .I5(\r9/t3/t0/p_0_in [2]),
        .O(\r9/p_0_out [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair340" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[2]_i_1__8 
       (.I0(\a10/k3a [2]),
        .I1(\a10/k4a [2]),
        .I2(\rf/p_0_in [2]),
        .O(\rf/p_4_out [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[30]_i_1 
       (.I0(\r1/t0/t1/p_1_in [6]),
        .I1(\r1/t0/t1/p_0_in [6]),
        .I2(\r1/t2/t3/p_0_in [6]),
        .I3(\r1/t1/t2/p_0_in [6]),
        .I4(k0b[30]),
        .I5(\r1/t3/t0/p_1_in [6]),
        .O(\r1/p_0_out [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[30]_i_1__0 
       (.I0(\r2/t0/t1/p_1_in [6]),
        .I1(\r2/t0/t1/p_0_in [6]),
        .I2(\r2/t2/t3/p_0_in [6]),
        .I3(\r2/t1/t2/p_0_in [6]),
        .I4(k1b[30]),
        .I5(\r2/t3/t0/p_1_in [6]),
        .O(\r2/p_0_out [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[30]_i_1__1 
       (.I0(\r3/t0/t1/p_1_in [6]),
        .I1(\r3/t0/t1/p_0_in [6]),
        .I2(\r3/t2/t3/p_0_in [6]),
        .I3(\r3/t1/t2/p_0_in [6]),
        .I4(k2b[30]),
        .I5(\r3/t3/t0/p_1_in [6]),
        .O(\r3/p_0_out [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[30]_i_1__2 
       (.I0(\r4/t0/t1/p_1_in [6]),
        .I1(\r4/t0/t1/p_0_in [6]),
        .I2(\r4/t2/t3/p_0_in [6]),
        .I3(\r4/t1/t2/p_0_in [6]),
        .I4(k3b[30]),
        .I5(\r4/t3/t0/p_1_in [6]),
        .O(\r4/p_0_out [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[30]_i_1__3 
       (.I0(\r5/t0/t1/p_1_in [6]),
        .I1(\r5/t0/t1/p_0_in [6]),
        .I2(\r5/t2/t3/p_0_in [6]),
        .I3(\r5/t1/t2/p_0_in [6]),
        .I4(k4b[30]),
        .I5(\r5/t3/t0/p_1_in [6]),
        .O(\r5/p_0_out [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[30]_i_1__4 
       (.I0(\r6/t0/t1/p_1_in [6]),
        .I1(\r6/t0/t1/p_0_in [6]),
        .I2(\r6/t2/t3/p_0_in [6]),
        .I3(\r6/t1/t2/p_0_in [6]),
        .I4(k5b[30]),
        .I5(\r6/t3/t0/p_1_in [6]),
        .O(\r6/p_0_out [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[30]_i_1__5 
       (.I0(\r7/t0/t1/p_1_in [6]),
        .I1(\r7/t0/t1/p_0_in [6]),
        .I2(\r7/t2/t3/p_0_in [6]),
        .I3(\r7/t1/t2/p_0_in [6]),
        .I4(k6b[30]),
        .I5(\r7/t3/t0/p_1_in [6]),
        .O(\r7/p_0_out [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[30]_i_1__6 
       (.I0(\r8/t0/t1/p_1_in [6]),
        .I1(\r8/t0/t1/p_0_in [6]),
        .I2(\r8/t2/t3/p_0_in [6]),
        .I3(\r8/t1/t2/p_0_in [6]),
        .I4(k7b[30]),
        .I5(\r8/t3/t0/p_1_in [6]),
        .O(\r8/p_0_out [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[30]_i_1__7 
       (.I0(\r9/t0/t1/p_1_in [6]),
        .I1(\r9/t0/t1/p_0_in [6]),
        .I2(\r9/t2/t3/p_0_in [6]),
        .I3(\r9/t1/t2/p_0_in [6]),
        .I4(k8b[30]),
        .I5(\r9/t3/t0/p_1_in [6]),
        .O(\r9/p_0_out [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair323" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[30]_i_1__8 
       (.I0(\a10/k3a [30]),
        .I1(\a10/k4a [30]),
        .I2(\rf/p_0_in [30]),
        .O(\rf/p_4_out [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[31]_i_1 
       (.I0(\r1/t0/t1/p_1_in [7]),
        .I1(\r1/t0/t1/p_0_in [7]),
        .I2(\r1/t2/t3/p_0_in [7]),
        .I3(\r1/t1/t2/p_0_in [7]),
        .I4(k0b[31]),
        .I5(\r1/t3/t0/p_1_in [7]),
        .O(\r1/p_0_out [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[31]_i_1__0 
       (.I0(\r2/t0/t1/p_1_in [7]),
        .I1(\r2/t0/t1/p_0_in [7]),
        .I2(\r2/t2/t3/p_0_in [7]),
        .I3(\r2/t1/t2/p_0_in [7]),
        .I4(k1b[31]),
        .I5(\r2/t3/t0/p_1_in [7]),
        .O(\r2/p_0_out [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[31]_i_1__1 
       (.I0(\r3/t0/t1/p_1_in [7]),
        .I1(\r3/t0/t1/p_0_in [7]),
        .I2(\r3/t2/t3/p_0_in [7]),
        .I3(\r3/t1/t2/p_0_in [7]),
        .I4(k2b[31]),
        .I5(\r3/t3/t0/p_1_in [7]),
        .O(\r3/p_0_out [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[31]_i_1__2 
       (.I0(\r4/t0/t1/p_1_in [7]),
        .I1(\r4/t0/t1/p_0_in [7]),
        .I2(\r4/t2/t3/p_0_in [7]),
        .I3(\r4/t1/t2/p_0_in [7]),
        .I4(k3b[31]),
        .I5(\r4/t3/t0/p_1_in [7]),
        .O(\r4/p_0_out [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[31]_i_1__3 
       (.I0(\r5/t0/t1/p_1_in [7]),
        .I1(\r5/t0/t1/p_0_in [7]),
        .I2(\r5/t2/t3/p_0_in [7]),
        .I3(\r5/t1/t2/p_0_in [7]),
        .I4(k4b[31]),
        .I5(\r5/t3/t0/p_1_in [7]),
        .O(\r5/p_0_out [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[31]_i_1__4 
       (.I0(\r6/t0/t1/p_1_in [7]),
        .I1(\r6/t0/t1/p_0_in [7]),
        .I2(\r6/t2/t3/p_0_in [7]),
        .I3(\r6/t1/t2/p_0_in [7]),
        .I4(k5b[31]),
        .I5(\r6/t3/t0/p_1_in [7]),
        .O(\r6/p_0_out [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[31]_i_1__5 
       (.I0(\r7/t0/t1/p_1_in [7]),
        .I1(\r7/t0/t1/p_0_in [7]),
        .I2(\r7/t2/t3/p_0_in [7]),
        .I3(\r7/t1/t2/p_0_in [7]),
        .I4(k6b[31]),
        .I5(\r7/t3/t0/p_1_in [7]),
        .O(\r7/p_0_out [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[31]_i_1__6 
       (.I0(\r8/t0/t1/p_1_in [7]),
        .I1(\r8/t0/t1/p_0_in [7]),
        .I2(\r8/t2/t3/p_0_in [7]),
        .I3(\r8/t1/t2/p_0_in [7]),
        .I4(k7b[31]),
        .I5(\r8/t3/t0/p_1_in [7]),
        .O(\r8/p_0_out [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[31]_i_1__7 
       (.I0(\r9/t0/t1/p_1_in [7]),
        .I1(\r9/t0/t1/p_0_in [7]),
        .I2(\r9/t2/t3/p_0_in [7]),
        .I3(\r9/t1/t2/p_0_in [7]),
        .I4(k8b[31]),
        .I5(\r9/t3/t0/p_1_in [7]),
        .O(\r9/p_0_out [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair324" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[31]_i_1__8 
       (.I0(\a10/k3a [31]),
        .I1(\a10/k4a [31]),
        .I2(\rf/p_0_in [31]),
        .O(\rf/p_4_out [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[32]_i_1 
       (.I0(\r1/t0/t2/p_0_in [0]),
        .I1(\r1/t2/t0/p_1_in [0]),
        .I2(\r1/t2/t0/p_0_in [0]),
        .I3(\r1/t1/t3/p_1_in [0]),
        .I4(k0b[32]),
        .I5(\r1/t3/t1/p_0_in [0]),
        .O(\r1/p_0_out [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[32]_i_1__0 
       (.I0(\r2/t0/t2/p_0_in [0]),
        .I1(\r2/t2/t0/p_1_in [0]),
        .I2(\r2/t2/t0/p_0_in [0]),
        .I3(\r2/t1/t3/p_1_in [0]),
        .I4(k1b[32]),
        .I5(\r2/t3/t1/p_0_in [0]),
        .O(\r2/p_0_out [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[32]_i_1__1 
       (.I0(\r3/t0/t2/p_0_in [0]),
        .I1(\r3/t2/t0/p_1_in [0]),
        .I2(\r3/t2/t0/p_0_in [0]),
        .I3(\r3/t1/t3/p_1_in [0]),
        .I4(k2b[32]),
        .I5(\r3/t3/t1/p_0_in [0]),
        .O(\r3/p_0_out [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[32]_i_1__2 
       (.I0(\r4/t0/t2/p_0_in [0]),
        .I1(\r4/t2/t0/p_1_in [0]),
        .I2(\r4/t2/t0/p_0_in [0]),
        .I3(\r4/t1/t3/p_1_in [0]),
        .I4(k3b[32]),
        .I5(\r4/t3/t1/p_0_in [0]),
        .O(\r4/p_0_out [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[32]_i_1__3 
       (.I0(\r5/t0/t2/p_0_in [0]),
        .I1(\r5/t2/t0/p_1_in [0]),
        .I2(\r5/t2/t0/p_0_in [0]),
        .I3(\r5/t1/t3/p_1_in [0]),
        .I4(k4b[32]),
        .I5(\r5/t3/t1/p_0_in [0]),
        .O(\r5/p_0_out [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[32]_i_1__4 
       (.I0(\r6/t0/t2/p_0_in [0]),
        .I1(\r6/t2/t0/p_1_in [0]),
        .I2(\r6/t2/t0/p_0_in [0]),
        .I3(\r6/t1/t3/p_1_in [0]),
        .I4(k5b[32]),
        .I5(\r6/t3/t1/p_0_in [0]),
        .O(\r6/p_0_out [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[32]_i_1__5 
       (.I0(\r7/t0/t2/p_0_in [0]),
        .I1(\r7/t2/t0/p_1_in [0]),
        .I2(\r7/t2/t0/p_0_in [0]),
        .I3(\r7/t1/t3/p_1_in [0]),
        .I4(k6b[32]),
        .I5(\r7/t3/t1/p_0_in [0]),
        .O(\r7/p_0_out [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[32]_i_1__6 
       (.I0(\r8/t0/t2/p_0_in [0]),
        .I1(\r8/t2/t0/p_1_in [0]),
        .I2(\r8/t2/t0/p_0_in [0]),
        .I3(\r8/t1/t3/p_1_in [0]),
        .I4(k7b[32]),
        .I5(\r8/t3/t1/p_0_in [0]),
        .O(\r8/p_0_out [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[32]_i_1__7 
       (.I0(\r9/t0/t2/p_0_in [0]),
        .I1(\r9/t2/t0/p_1_in [0]),
        .I2(\r9/t2/t0/p_0_in [0]),
        .I3(\r9/t1/t3/p_1_in [0]),
        .I4(k8b[32]),
        .I5(\r9/t3/t1/p_0_in [0]),
        .O(\r9/p_0_out [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair374" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[32]_i_1__8 
       (.I0(\a10/k2a [0]),
        .I1(\a10/k4a [0]),
        .I2(\rf/p_1_in [0]),
        .O(\rf/p_4_out [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[33]_i_1 
       (.I0(\r1/t0/t2/p_0_in [1]),
        .I1(\r1/t2/t0/p_1_in [1]),
        .I2(\r1/t2/t0/p_0_in [1]),
        .I3(\r1/t1/t3/p_1_in [1]),
        .I4(k0b[33]),
        .I5(\r1/t3/t1/p_0_in [1]),
        .O(\r1/p_0_out [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[33]_i_1__0 
       (.I0(\r2/t0/t2/p_0_in [1]),
        .I1(\r2/t2/t0/p_1_in [1]),
        .I2(\r2/t2/t0/p_0_in [1]),
        .I3(\r2/t1/t3/p_1_in [1]),
        .I4(k1b[33]),
        .I5(\r2/t3/t1/p_0_in [1]),
        .O(\r2/p_0_out [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[33]_i_1__1 
       (.I0(\r3/t0/t2/p_0_in [1]),
        .I1(\r3/t2/t0/p_1_in [1]),
        .I2(\r3/t2/t0/p_0_in [1]),
        .I3(\r3/t1/t3/p_1_in [1]),
        .I4(k2b[33]),
        .I5(\r3/t3/t1/p_0_in [1]),
        .O(\r3/p_0_out [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[33]_i_1__2 
       (.I0(\r4/t0/t2/p_0_in [1]),
        .I1(\r4/t2/t0/p_1_in [1]),
        .I2(\r4/t2/t0/p_0_in [1]),
        .I3(\r4/t1/t3/p_1_in [1]),
        .I4(k3b[33]),
        .I5(\r4/t3/t1/p_0_in [1]),
        .O(\r4/p_0_out [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[33]_i_1__3 
       (.I0(\r5/t0/t2/p_0_in [1]),
        .I1(\r5/t2/t0/p_1_in [1]),
        .I2(\r5/t2/t0/p_0_in [1]),
        .I3(\r5/t1/t3/p_1_in [1]),
        .I4(k4b[33]),
        .I5(\r5/t3/t1/p_0_in [1]),
        .O(\r5/p_0_out [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[33]_i_1__4 
       (.I0(\r6/t0/t2/p_0_in [1]),
        .I1(\r6/t2/t0/p_1_in [1]),
        .I2(\r6/t2/t0/p_0_in [1]),
        .I3(\r6/t1/t3/p_1_in [1]),
        .I4(k5b[33]),
        .I5(\r6/t3/t1/p_0_in [1]),
        .O(\r6/p_0_out [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[33]_i_1__5 
       (.I0(\r7/t0/t2/p_0_in [1]),
        .I1(\r7/t2/t0/p_1_in [1]),
        .I2(\r7/t2/t0/p_0_in [1]),
        .I3(\r7/t1/t3/p_1_in [1]),
        .I4(k6b[33]),
        .I5(\r7/t3/t1/p_0_in [1]),
        .O(\r7/p_0_out [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[33]_i_1__6 
       (.I0(\r8/t0/t2/p_0_in [1]),
        .I1(\r8/t2/t0/p_1_in [1]),
        .I2(\r8/t2/t0/p_0_in [1]),
        .I3(\r8/t1/t3/p_1_in [1]),
        .I4(k7b[33]),
        .I5(\r8/t3/t1/p_0_in [1]),
        .O(\r8/p_0_out [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[33]_i_1__7 
       (.I0(\r9/t0/t2/p_0_in [1]),
        .I1(\r9/t2/t0/p_1_in [1]),
        .I2(\r9/t2/t0/p_0_in [1]),
        .I3(\r9/t1/t3/p_1_in [1]),
        .I4(k8b[33]),
        .I5(\r9/t3/t1/p_0_in [1]),
        .O(\r9/p_0_out [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair373" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[33]_i_1__8 
       (.I0(\a10/k2a [1]),
        .I1(\a10/k4a [1]),
        .I2(\rf/p_1_in [1]),
        .O(\rf/p_4_out [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[34]_i_1 
       (.I0(\r1/t0/t2/p_0_in [2]),
        .I1(\r1/t2/t0/p_1_in [2]),
        .I2(\r1/t2/t0/p_0_in [2]),
        .I3(\r1/t1/t3/p_1_in [2]),
        .I4(k0b[34]),
        .I5(\r1/t3/t1/p_0_in [2]),
        .O(\r1/p_0_out [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[34]_i_1__0 
       (.I0(\r2/t0/t2/p_0_in [2]),
        .I1(\r2/t2/t0/p_1_in [2]),
        .I2(\r2/t2/t0/p_0_in [2]),
        .I3(\r2/t1/t3/p_1_in [2]),
        .I4(k1b[34]),
        .I5(\r2/t3/t1/p_0_in [2]),
        .O(\r2/p_0_out [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[34]_i_1__1 
       (.I0(\r3/t0/t2/p_0_in [2]),
        .I1(\r3/t2/t0/p_1_in [2]),
        .I2(\r3/t2/t0/p_0_in [2]),
        .I3(\r3/t1/t3/p_1_in [2]),
        .I4(k2b[34]),
        .I5(\r3/t3/t1/p_0_in [2]),
        .O(\r3/p_0_out [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[34]_i_1__2 
       (.I0(\r4/t0/t2/p_0_in [2]),
        .I1(\r4/t2/t0/p_1_in [2]),
        .I2(\r4/t2/t0/p_0_in [2]),
        .I3(\r4/t1/t3/p_1_in [2]),
        .I4(k3b[34]),
        .I5(\r4/t3/t1/p_0_in [2]),
        .O(\r4/p_0_out [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[34]_i_1__3 
       (.I0(\r5/t0/t2/p_0_in [2]),
        .I1(\r5/t2/t0/p_1_in [2]),
        .I2(\r5/t2/t0/p_0_in [2]),
        .I3(\r5/t1/t3/p_1_in [2]),
        .I4(k4b[34]),
        .I5(\r5/t3/t1/p_0_in [2]),
        .O(\r5/p_0_out [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[34]_i_1__4 
       (.I0(\r6/t0/t2/p_0_in [2]),
        .I1(\r6/t2/t0/p_1_in [2]),
        .I2(\r6/t2/t0/p_0_in [2]),
        .I3(\r6/t1/t3/p_1_in [2]),
        .I4(k5b[34]),
        .I5(\r6/t3/t1/p_0_in [2]),
        .O(\r6/p_0_out [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[34]_i_1__5 
       (.I0(\r7/t0/t2/p_0_in [2]),
        .I1(\r7/t2/t0/p_1_in [2]),
        .I2(\r7/t2/t0/p_0_in [2]),
        .I3(\r7/t1/t3/p_1_in [2]),
        .I4(k6b[34]),
        .I5(\r7/t3/t1/p_0_in [2]),
        .O(\r7/p_0_out [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[34]_i_1__6 
       (.I0(\r8/t0/t2/p_0_in [2]),
        .I1(\r8/t2/t0/p_1_in [2]),
        .I2(\r8/t2/t0/p_0_in [2]),
        .I3(\r8/t1/t3/p_1_in [2]),
        .I4(k7b[34]),
        .I5(\r8/t3/t1/p_0_in [2]),
        .O(\r8/p_0_out [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[34]_i_1__7 
       (.I0(\r9/t0/t2/p_0_in [2]),
        .I1(\r9/t2/t0/p_1_in [2]),
        .I2(\r9/t2/t0/p_0_in [2]),
        .I3(\r9/t1/t3/p_1_in [2]),
        .I4(k8b[34]),
        .I5(\r9/t3/t1/p_0_in [2]),
        .O(\r9/p_0_out [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair372" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[34]_i_1__8 
       (.I0(\a10/k2a [2]),
        .I1(\a10/k4a [2]),
        .I2(\rf/p_1_in [2]),
        .O(\rf/p_4_out [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[35]_i_1 
       (.I0(\r1/t0/t2/p_0_in [3]),
        .I1(\r1/t2/t0/p_1_in [3]),
        .I2(\r1/t2/t0/p_0_in [3]),
        .I3(\r1/t1/t3/p_1_in [3]),
        .I4(k0b[35]),
        .I5(\r1/t3/t1/p_0_in [3]),
        .O(\r1/p_0_out [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[35]_i_1__0 
       (.I0(\r2/t0/t2/p_0_in [3]),
        .I1(\r2/t2/t0/p_1_in [3]),
        .I2(\r2/t2/t0/p_0_in [3]),
        .I3(\r2/t1/t3/p_1_in [3]),
        .I4(k1b[35]),
        .I5(\r2/t3/t1/p_0_in [3]),
        .O(\r2/p_0_out [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[35]_i_1__1 
       (.I0(\r3/t0/t2/p_0_in [3]),
        .I1(\r3/t2/t0/p_1_in [3]),
        .I2(\r3/t2/t0/p_0_in [3]),
        .I3(\r3/t1/t3/p_1_in [3]),
        .I4(k2b[35]),
        .I5(\r3/t3/t1/p_0_in [3]),
        .O(\r3/p_0_out [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[35]_i_1__2 
       (.I0(\r4/t0/t2/p_0_in [3]),
        .I1(\r4/t2/t0/p_1_in [3]),
        .I2(\r4/t2/t0/p_0_in [3]),
        .I3(\r4/t1/t3/p_1_in [3]),
        .I4(k3b[35]),
        .I5(\r4/t3/t1/p_0_in [3]),
        .O(\r4/p_0_out [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[35]_i_1__3 
       (.I0(\r5/t0/t2/p_0_in [3]),
        .I1(\r5/t2/t0/p_1_in [3]),
        .I2(\r5/t2/t0/p_0_in [3]),
        .I3(\r5/t1/t3/p_1_in [3]),
        .I4(k4b[35]),
        .I5(\r5/t3/t1/p_0_in [3]),
        .O(\r5/p_0_out [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[35]_i_1__4 
       (.I0(\r6/t0/t2/p_0_in [3]),
        .I1(\r6/t2/t0/p_1_in [3]),
        .I2(\r6/t2/t0/p_0_in [3]),
        .I3(\r6/t1/t3/p_1_in [3]),
        .I4(k5b[35]),
        .I5(\r6/t3/t1/p_0_in [3]),
        .O(\r6/p_0_out [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[35]_i_1__5 
       (.I0(\r7/t0/t2/p_0_in [3]),
        .I1(\r7/t2/t0/p_1_in [3]),
        .I2(\r7/t2/t0/p_0_in [3]),
        .I3(\r7/t1/t3/p_1_in [3]),
        .I4(k6b[35]),
        .I5(\r7/t3/t1/p_0_in [3]),
        .O(\r7/p_0_out [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[35]_i_1__6 
       (.I0(\r8/t0/t2/p_0_in [3]),
        .I1(\r8/t2/t0/p_1_in [3]),
        .I2(\r8/t2/t0/p_0_in [3]),
        .I3(\r8/t1/t3/p_1_in [3]),
        .I4(k7b[35]),
        .I5(\r8/t3/t1/p_0_in [3]),
        .O(\r8/p_0_out [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[35]_i_1__7 
       (.I0(\r9/t0/t2/p_0_in [3]),
        .I1(\r9/t2/t0/p_1_in [3]),
        .I2(\r9/t2/t0/p_0_in [3]),
        .I3(\r9/t1/t3/p_1_in [3]),
        .I4(k8b[35]),
        .I5(\r9/t3/t1/p_0_in [3]),
        .O(\r9/p_0_out [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair371" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[35]_i_1__8 
       (.I0(\a10/k2a [3]),
        .I1(\a10/k4a [3]),
        .I2(\rf/p_1_in [3]),
        .O(\rf/p_4_out [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[36]_i_1 
       (.I0(\r1/t0/t2/p_0_in [4]),
        .I1(\r1/t2/t0/p_1_in [4]),
        .I2(\r1/t2/t0/p_0_in [4]),
        .I3(\r1/t1/t3/p_1_in [4]),
        .I4(k0b[36]),
        .I5(\r1/t3/t1/p_0_in [4]),
        .O(\r1/p_0_out [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[36]_i_1__0 
       (.I0(\r2/t0/t2/p_0_in [4]),
        .I1(\r2/t2/t0/p_1_in [4]),
        .I2(\r2/t2/t0/p_0_in [4]),
        .I3(\r2/t1/t3/p_1_in [4]),
        .I4(k1b[36]),
        .I5(\r2/t3/t1/p_0_in [4]),
        .O(\r2/p_0_out [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[36]_i_1__1 
       (.I0(\r3/t0/t2/p_0_in [4]),
        .I1(\r3/t2/t0/p_1_in [4]),
        .I2(\r3/t2/t0/p_0_in [4]),
        .I3(\r3/t1/t3/p_1_in [4]),
        .I4(k2b[36]),
        .I5(\r3/t3/t1/p_0_in [4]),
        .O(\r3/p_0_out [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[36]_i_1__2 
       (.I0(\r4/t0/t2/p_0_in [4]),
        .I1(\r4/t2/t0/p_1_in [4]),
        .I2(\r4/t2/t0/p_0_in [4]),
        .I3(\r4/t1/t3/p_1_in [4]),
        .I4(k3b[36]),
        .I5(\r4/t3/t1/p_0_in [4]),
        .O(\r4/p_0_out [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[36]_i_1__3 
       (.I0(\r5/t0/t2/p_0_in [4]),
        .I1(\r5/t2/t0/p_1_in [4]),
        .I2(\r5/t2/t0/p_0_in [4]),
        .I3(\r5/t1/t3/p_1_in [4]),
        .I4(k4b[36]),
        .I5(\r5/t3/t1/p_0_in [4]),
        .O(\r5/p_0_out [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[36]_i_1__4 
       (.I0(\r6/t0/t2/p_0_in [4]),
        .I1(\r6/t2/t0/p_1_in [4]),
        .I2(\r6/t2/t0/p_0_in [4]),
        .I3(\r6/t1/t3/p_1_in [4]),
        .I4(k5b[36]),
        .I5(\r6/t3/t1/p_0_in [4]),
        .O(\r6/p_0_out [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[36]_i_1__5 
       (.I0(\r7/t0/t2/p_0_in [4]),
        .I1(\r7/t2/t0/p_1_in [4]),
        .I2(\r7/t2/t0/p_0_in [4]),
        .I3(\r7/t1/t3/p_1_in [4]),
        .I4(k6b[36]),
        .I5(\r7/t3/t1/p_0_in [4]),
        .O(\r7/p_0_out [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[36]_i_1__6 
       (.I0(\r8/t0/t2/p_0_in [4]),
        .I1(\r8/t2/t0/p_1_in [4]),
        .I2(\r8/t2/t0/p_0_in [4]),
        .I3(\r8/t1/t3/p_1_in [4]),
        .I4(k7b[36]),
        .I5(\r8/t3/t1/p_0_in [4]),
        .O(\r8/p_0_out [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[36]_i_1__7 
       (.I0(\r9/t0/t2/p_0_in [4]),
        .I1(\r9/t2/t0/p_1_in [4]),
        .I2(\r9/t2/t0/p_0_in [4]),
        .I3(\r9/t1/t3/p_1_in [4]),
        .I4(k8b[36]),
        .I5(\r9/t3/t1/p_0_in [4]),
        .O(\r9/p_0_out [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair370" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[36]_i_1__8 
       (.I0(\a10/k2a [4]),
        .I1(\a10/k4a [4]),
        .I2(\rf/p_1_in [4]),
        .O(\rf/p_4_out [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[37]_i_1 
       (.I0(\r1/t0/t2/p_0_in [5]),
        .I1(\r1/t2/t0/p_1_in [5]),
        .I2(\r1/t2/t0/p_0_in [5]),
        .I3(\r1/t1/t3/p_1_in [5]),
        .I4(k0b[37]),
        .I5(\r1/t3/t1/p_0_in [5]),
        .O(\r1/p_0_out [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[37]_i_1__0 
       (.I0(\r2/t0/t2/p_0_in [5]),
        .I1(\r2/t2/t0/p_1_in [5]),
        .I2(\r2/t2/t0/p_0_in [5]),
        .I3(\r2/t1/t3/p_1_in [5]),
        .I4(k1b[37]),
        .I5(\r2/t3/t1/p_0_in [5]),
        .O(\r2/p_0_out [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[37]_i_1__1 
       (.I0(\r3/t0/t2/p_0_in [5]),
        .I1(\r3/t2/t0/p_1_in [5]),
        .I2(\r3/t2/t0/p_0_in [5]),
        .I3(\r3/t1/t3/p_1_in [5]),
        .I4(k2b[37]),
        .I5(\r3/t3/t1/p_0_in [5]),
        .O(\r3/p_0_out [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[37]_i_1__2 
       (.I0(\r4/t0/t2/p_0_in [5]),
        .I1(\r4/t2/t0/p_1_in [5]),
        .I2(\r4/t2/t0/p_0_in [5]),
        .I3(\r4/t1/t3/p_1_in [5]),
        .I4(k3b[37]),
        .I5(\r4/t3/t1/p_0_in [5]),
        .O(\r4/p_0_out [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[37]_i_1__3 
       (.I0(\r5/t0/t2/p_0_in [5]),
        .I1(\r5/t2/t0/p_1_in [5]),
        .I2(\r5/t2/t0/p_0_in [5]),
        .I3(\r5/t1/t3/p_1_in [5]),
        .I4(k4b[37]),
        .I5(\r5/t3/t1/p_0_in [5]),
        .O(\r5/p_0_out [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[37]_i_1__4 
       (.I0(\r6/t0/t2/p_0_in [5]),
        .I1(\r6/t2/t0/p_1_in [5]),
        .I2(\r6/t2/t0/p_0_in [5]),
        .I3(\r6/t1/t3/p_1_in [5]),
        .I4(k5b[37]),
        .I5(\r6/t3/t1/p_0_in [5]),
        .O(\r6/p_0_out [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[37]_i_1__5 
       (.I0(\r7/t0/t2/p_0_in [5]),
        .I1(\r7/t2/t0/p_1_in [5]),
        .I2(\r7/t2/t0/p_0_in [5]),
        .I3(\r7/t1/t3/p_1_in [5]),
        .I4(k6b[37]),
        .I5(\r7/t3/t1/p_0_in [5]),
        .O(\r7/p_0_out [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[37]_i_1__6 
       (.I0(\r8/t0/t2/p_0_in [5]),
        .I1(\r8/t2/t0/p_1_in [5]),
        .I2(\r8/t2/t0/p_0_in [5]),
        .I3(\r8/t1/t3/p_1_in [5]),
        .I4(k7b[37]),
        .I5(\r8/t3/t1/p_0_in [5]),
        .O(\r8/p_0_out [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[37]_i_1__7 
       (.I0(\r9/t0/t2/p_0_in [5]),
        .I1(\r9/t2/t0/p_1_in [5]),
        .I2(\r9/t2/t0/p_0_in [5]),
        .I3(\r9/t1/t3/p_1_in [5]),
        .I4(k8b[37]),
        .I5(\r9/t3/t1/p_0_in [5]),
        .O(\r9/p_0_out [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair369" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[37]_i_1__8 
       (.I0(\a10/k2a [5]),
        .I1(\a10/k4a [5]),
        .I2(\rf/p_1_in [5]),
        .O(\rf/p_4_out [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[38]_i_1 
       (.I0(\r1/t0/t2/p_0_in [6]),
        .I1(\r1/t2/t0/p_1_in [6]),
        .I2(\r1/t2/t0/p_0_in [6]),
        .I3(\r1/t1/t3/p_1_in [6]),
        .I4(k0b[38]),
        .I5(\r1/t3/t1/p_0_in [6]),
        .O(\r1/p_0_out [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[38]_i_1__0 
       (.I0(\r2/t0/t2/p_0_in [6]),
        .I1(\r2/t2/t0/p_1_in [6]),
        .I2(\r2/t2/t0/p_0_in [6]),
        .I3(\r2/t1/t3/p_1_in [6]),
        .I4(k1b[38]),
        .I5(\r2/t3/t1/p_0_in [6]),
        .O(\r2/p_0_out [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[38]_i_1__1 
       (.I0(\r3/t0/t2/p_0_in [6]),
        .I1(\r3/t2/t0/p_1_in [6]),
        .I2(\r3/t2/t0/p_0_in [6]),
        .I3(\r3/t1/t3/p_1_in [6]),
        .I4(k2b[38]),
        .I5(\r3/t3/t1/p_0_in [6]),
        .O(\r3/p_0_out [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[38]_i_1__2 
       (.I0(\r4/t0/t2/p_0_in [6]),
        .I1(\r4/t2/t0/p_1_in [6]),
        .I2(\r4/t2/t0/p_0_in [6]),
        .I3(\r4/t1/t3/p_1_in [6]),
        .I4(k3b[38]),
        .I5(\r4/t3/t1/p_0_in [6]),
        .O(\r4/p_0_out [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[38]_i_1__3 
       (.I0(\r5/t0/t2/p_0_in [6]),
        .I1(\r5/t2/t0/p_1_in [6]),
        .I2(\r5/t2/t0/p_0_in [6]),
        .I3(\r5/t1/t3/p_1_in [6]),
        .I4(k4b[38]),
        .I5(\r5/t3/t1/p_0_in [6]),
        .O(\r5/p_0_out [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[38]_i_1__4 
       (.I0(\r6/t0/t2/p_0_in [6]),
        .I1(\r6/t2/t0/p_1_in [6]),
        .I2(\r6/t2/t0/p_0_in [6]),
        .I3(\r6/t1/t3/p_1_in [6]),
        .I4(k5b[38]),
        .I5(\r6/t3/t1/p_0_in [6]),
        .O(\r6/p_0_out [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[38]_i_1__5 
       (.I0(\r7/t0/t2/p_0_in [6]),
        .I1(\r7/t2/t0/p_1_in [6]),
        .I2(\r7/t2/t0/p_0_in [6]),
        .I3(\r7/t1/t3/p_1_in [6]),
        .I4(k6b[38]),
        .I5(\r7/t3/t1/p_0_in [6]),
        .O(\r7/p_0_out [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[38]_i_1__6 
       (.I0(\r8/t0/t2/p_0_in [6]),
        .I1(\r8/t2/t0/p_1_in [6]),
        .I2(\r8/t2/t0/p_0_in [6]),
        .I3(\r8/t1/t3/p_1_in [6]),
        .I4(k7b[38]),
        .I5(\r8/t3/t1/p_0_in [6]),
        .O(\r8/p_0_out [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[38]_i_1__7 
       (.I0(\r9/t0/t2/p_0_in [6]),
        .I1(\r9/t2/t0/p_1_in [6]),
        .I2(\r9/t2/t0/p_0_in [6]),
        .I3(\r9/t1/t3/p_1_in [6]),
        .I4(k8b[38]),
        .I5(\r9/t3/t1/p_0_in [6]),
        .O(\r9/p_0_out [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair368" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[38]_i_1__8 
       (.I0(\a10/k2a [6]),
        .I1(\a10/k4a [6]),
        .I2(\rf/p_1_in [6]),
        .O(\rf/p_4_out [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[39]_i_1 
       (.I0(\r1/t0/t2/p_0_in [7]),
        .I1(\r1/t2/t0/p_1_in [7]),
        .I2(\r1/t2/t0/p_0_in [7]),
        .I3(\r1/t1/t3/p_1_in [7]),
        .I4(k0b[39]),
        .I5(\r1/t3/t1/p_0_in [7]),
        .O(\r1/p_0_out [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[39]_i_1__0 
       (.I0(\r2/t0/t2/p_0_in [7]),
        .I1(\r2/t2/t0/p_1_in [7]),
        .I2(\r2/t2/t0/p_0_in [7]),
        .I3(\r2/t1/t3/p_1_in [7]),
        .I4(k1b[39]),
        .I5(\r2/t3/t1/p_0_in [7]),
        .O(\r2/p_0_out [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[39]_i_1__1 
       (.I0(\r3/t0/t2/p_0_in [7]),
        .I1(\r3/t2/t0/p_1_in [7]),
        .I2(\r3/t2/t0/p_0_in [7]),
        .I3(\r3/t1/t3/p_1_in [7]),
        .I4(k2b[39]),
        .I5(\r3/t3/t1/p_0_in [7]),
        .O(\r3/p_0_out [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[39]_i_1__2 
       (.I0(\r4/t0/t2/p_0_in [7]),
        .I1(\r4/t2/t0/p_1_in [7]),
        .I2(\r4/t2/t0/p_0_in [7]),
        .I3(\r4/t1/t3/p_1_in [7]),
        .I4(k3b[39]),
        .I5(\r4/t3/t1/p_0_in [7]),
        .O(\r4/p_0_out [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[39]_i_1__3 
       (.I0(\r5/t0/t2/p_0_in [7]),
        .I1(\r5/t2/t0/p_1_in [7]),
        .I2(\r5/t2/t0/p_0_in [7]),
        .I3(\r5/t1/t3/p_1_in [7]),
        .I4(k4b[39]),
        .I5(\r5/t3/t1/p_0_in [7]),
        .O(\r5/p_0_out [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[39]_i_1__4 
       (.I0(\r6/t0/t2/p_0_in [7]),
        .I1(\r6/t2/t0/p_1_in [7]),
        .I2(\r6/t2/t0/p_0_in [7]),
        .I3(\r6/t1/t3/p_1_in [7]),
        .I4(k5b[39]),
        .I5(\r6/t3/t1/p_0_in [7]),
        .O(\r6/p_0_out [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[39]_i_1__5 
       (.I0(\r7/t0/t2/p_0_in [7]),
        .I1(\r7/t2/t0/p_1_in [7]),
        .I2(\r7/t2/t0/p_0_in [7]),
        .I3(\r7/t1/t3/p_1_in [7]),
        .I4(k6b[39]),
        .I5(\r7/t3/t1/p_0_in [7]),
        .O(\r7/p_0_out [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[39]_i_1__6 
       (.I0(\r8/t0/t2/p_0_in [7]),
        .I1(\r8/t2/t0/p_1_in [7]),
        .I2(\r8/t2/t0/p_0_in [7]),
        .I3(\r8/t1/t3/p_1_in [7]),
        .I4(k7b[39]),
        .I5(\r8/t3/t1/p_0_in [7]),
        .O(\r8/p_0_out [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[39]_i_1__7 
       (.I0(\r9/t0/t2/p_0_in [7]),
        .I1(\r9/t2/t0/p_1_in [7]),
        .I2(\r9/t2/t0/p_0_in [7]),
        .I3(\r9/t1/t3/p_1_in [7]),
        .I4(k8b[39]),
        .I5(\r9/t3/t1/p_0_in [7]),
        .O(\r9/p_0_out [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair367" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[39]_i_1__8 
       (.I0(\a10/k2a [7]),
        .I1(\a10/k4a [7]),
        .I2(\rf/p_1_in [7]),
        .O(\rf/p_4_out [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[3]_i_1 
       (.I0(\r1/t0/t1/p_0_in [3]),
        .I1(\r1/t2/t3/p_1_in [3]),
        .I2(\r1/t1/t2/p_0_in [3]),
        .I3(k0b[3]),
        .I4(\r1/t3/t0/p_1_in [3]),
        .I5(\r1/t3/t0/p_0_in [3]),
        .O(\r1/p_0_out [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[3]_i_1__0 
       (.I0(\r2/t0/t1/p_0_in [3]),
        .I1(\r2/t2/t3/p_1_in [3]),
        .I2(\r2/t1/t2/p_0_in [3]),
        .I3(k1b[3]),
        .I4(\r2/t3/t0/p_1_in [3]),
        .I5(\r2/t3/t0/p_0_in [3]),
        .O(\r2/p_0_out [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[3]_i_1__1 
       (.I0(\r3/t0/t1/p_0_in [3]),
        .I1(\r3/t2/t3/p_1_in [3]),
        .I2(\r3/t1/t2/p_0_in [3]),
        .I3(k2b[3]),
        .I4(\r3/t3/t0/p_1_in [3]),
        .I5(\r3/t3/t0/p_0_in [3]),
        .O(\r3/p_0_out [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[3]_i_1__2 
       (.I0(\r4/t0/t1/p_0_in [3]),
        .I1(\r4/t2/t3/p_1_in [3]),
        .I2(\r4/t1/t2/p_0_in [3]),
        .I3(k3b[3]),
        .I4(\r4/t3/t0/p_1_in [3]),
        .I5(\r4/t3/t0/p_0_in [3]),
        .O(\r4/p_0_out [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[3]_i_1__3 
       (.I0(\r5/t0/t1/p_0_in [3]),
        .I1(\r5/t2/t3/p_1_in [3]),
        .I2(\r5/t1/t2/p_0_in [3]),
        .I3(k4b[3]),
        .I4(\r5/t3/t0/p_1_in [3]),
        .I5(\r5/t3/t0/p_0_in [3]),
        .O(\r5/p_0_out [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[3]_i_1__4 
       (.I0(\r6/t0/t1/p_0_in [3]),
        .I1(\r6/t2/t3/p_1_in [3]),
        .I2(\r6/t1/t2/p_0_in [3]),
        .I3(k5b[3]),
        .I4(\r6/t3/t0/p_1_in [3]),
        .I5(\r6/t3/t0/p_0_in [3]),
        .O(\r6/p_0_out [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[3]_i_1__5 
       (.I0(\r7/t0/t1/p_0_in [3]),
        .I1(\r7/t2/t3/p_1_in [3]),
        .I2(\r7/t1/t2/p_0_in [3]),
        .I3(k6b[3]),
        .I4(\r7/t3/t0/p_1_in [3]),
        .I5(\r7/t3/t0/p_0_in [3]),
        .O(\r7/p_0_out [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[3]_i_1__6 
       (.I0(\r8/t0/t1/p_0_in [3]),
        .I1(\r8/t2/t3/p_1_in [3]),
        .I2(\r8/t1/t2/p_0_in [3]),
        .I3(k7b[3]),
        .I4(\r8/t3/t0/p_1_in [3]),
        .I5(\r8/t3/t0/p_0_in [3]),
        .O(\r8/p_0_out [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[3]_i_1__7 
       (.I0(\r9/t0/t1/p_0_in [3]),
        .I1(\r9/t2/t3/p_1_in [3]),
        .I2(\r9/t1/t2/p_0_in [3]),
        .I3(k8b[3]),
        .I4(\r9/t3/t0/p_1_in [3]),
        .I5(\r9/t3/t0/p_0_in [3]),
        .O(\r9/p_0_out [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair339" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[3]_i_1__8 
       (.I0(\a10/k3a [3]),
        .I1(\a10/k4a [3]),
        .I2(\rf/p_0_in [3]),
        .O(\rf/p_4_out [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[40]_i_1 
       (.I0(\r1/t0/t2/p_1_in [0]),
        .I1(\r1/t2/t0/p_0_in [0]),
        .I2(\r1/t1/t3/p_1_in [0]),
        .I3(\r1/t1/t3/p_0_in [0]),
        .I4(k0b[40]),
        .I5(\r1/t3/t1/p_0_in [0]),
        .O(\r1/p_0_out [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[40]_i_1__0 
       (.I0(\r2/t0/t2/p_1_in [0]),
        .I1(\r2/t2/t0/p_0_in [0]),
        .I2(\r2/t1/t3/p_1_in [0]),
        .I3(\r2/t1/t3/p_0_in [0]),
        .I4(k1b[40]),
        .I5(\r2/t3/t1/p_0_in [0]),
        .O(\r2/p_0_out [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[40]_i_1__1 
       (.I0(\r3/t0/t2/p_1_in [0]),
        .I1(\r3/t2/t0/p_0_in [0]),
        .I2(\r3/t1/t3/p_1_in [0]),
        .I3(\r3/t1/t3/p_0_in [0]),
        .I4(k2b[40]),
        .I5(\r3/t3/t1/p_0_in [0]),
        .O(\r3/p_0_out [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[40]_i_1__2 
       (.I0(\r4/t0/t2/p_1_in [0]),
        .I1(\r4/t2/t0/p_0_in [0]),
        .I2(\r4/t1/t3/p_1_in [0]),
        .I3(\r4/t1/t3/p_0_in [0]),
        .I4(k3b[40]),
        .I5(\r4/t3/t1/p_0_in [0]),
        .O(\r4/p_0_out [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[40]_i_1__3 
       (.I0(\r5/t0/t2/p_1_in [0]),
        .I1(\r5/t2/t0/p_0_in [0]),
        .I2(\r5/t1/t3/p_1_in [0]),
        .I3(\r5/t1/t3/p_0_in [0]),
        .I4(k4b[40]),
        .I5(\r5/t3/t1/p_0_in [0]),
        .O(\r5/p_0_out [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[40]_i_1__4 
       (.I0(\r6/t0/t2/p_1_in [0]),
        .I1(\r6/t2/t0/p_0_in [0]),
        .I2(\r6/t1/t3/p_1_in [0]),
        .I3(\r6/t1/t3/p_0_in [0]),
        .I4(k5b[40]),
        .I5(\r6/t3/t1/p_0_in [0]),
        .O(\r6/p_0_out [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[40]_i_1__5 
       (.I0(\r7/t0/t2/p_1_in [0]),
        .I1(\r7/t2/t0/p_0_in [0]),
        .I2(\r7/t1/t3/p_1_in [0]),
        .I3(\r7/t1/t3/p_0_in [0]),
        .I4(k6b[40]),
        .I5(\r7/t3/t1/p_0_in [0]),
        .O(\r7/p_0_out [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[40]_i_1__6 
       (.I0(\r8/t0/t2/p_1_in [0]),
        .I1(\r8/t2/t0/p_0_in [0]),
        .I2(\r8/t1/t3/p_1_in [0]),
        .I3(\r8/t1/t3/p_0_in [0]),
        .I4(k7b[40]),
        .I5(\r8/t3/t1/p_0_in [0]),
        .O(\r8/p_0_out [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[40]_i_1__7 
       (.I0(\r9/t0/t2/p_1_in [0]),
        .I1(\r9/t2/t0/p_0_in [0]),
        .I2(\r9/t1/t3/p_1_in [0]),
        .I3(\r9/t1/t3/p_0_in [0]),
        .I4(k8b[40]),
        .I5(\r9/t3/t1/p_0_in [0]),
        .O(\r9/p_0_out [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair366" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[40]_i_1__8 
       (.I0(\a10/k2a [8]),
        .I1(\a10/k4a [8]),
        .I2(\rf/p_1_in [8]),
        .O(\rf/p_4_out [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[41]_i_1 
       (.I0(\r1/t0/t2/p_1_in [1]),
        .I1(\r1/t2/t0/p_0_in [1]),
        .I2(\r1/t1/t3/p_1_in [1]),
        .I3(\r1/t1/t3/p_0_in [1]),
        .I4(k0b[41]),
        .I5(\r1/t3/t1/p_0_in [1]),
        .O(\r1/p_0_out [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[41]_i_1__0 
       (.I0(\r2/t0/t2/p_1_in [1]),
        .I1(\r2/t2/t0/p_0_in [1]),
        .I2(\r2/t1/t3/p_1_in [1]),
        .I3(\r2/t1/t3/p_0_in [1]),
        .I4(k1b[41]),
        .I5(\r2/t3/t1/p_0_in [1]),
        .O(\r2/p_0_out [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[41]_i_1__1 
       (.I0(\r3/t0/t2/p_1_in [1]),
        .I1(\r3/t2/t0/p_0_in [1]),
        .I2(\r3/t1/t3/p_1_in [1]),
        .I3(\r3/t1/t3/p_0_in [1]),
        .I4(k2b[41]),
        .I5(\r3/t3/t1/p_0_in [1]),
        .O(\r3/p_0_out [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[41]_i_1__2 
       (.I0(\r4/t0/t2/p_1_in [1]),
        .I1(\r4/t2/t0/p_0_in [1]),
        .I2(\r4/t1/t3/p_1_in [1]),
        .I3(\r4/t1/t3/p_0_in [1]),
        .I4(k3b[41]),
        .I5(\r4/t3/t1/p_0_in [1]),
        .O(\r4/p_0_out [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[41]_i_1__3 
       (.I0(\r5/t0/t2/p_1_in [1]),
        .I1(\r5/t2/t0/p_0_in [1]),
        .I2(\r5/t1/t3/p_1_in [1]),
        .I3(\r5/t1/t3/p_0_in [1]),
        .I4(k4b[41]),
        .I5(\r5/t3/t1/p_0_in [1]),
        .O(\r5/p_0_out [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[41]_i_1__4 
       (.I0(\r6/t0/t2/p_1_in [1]),
        .I1(\r6/t2/t0/p_0_in [1]),
        .I2(\r6/t1/t3/p_1_in [1]),
        .I3(\r6/t1/t3/p_0_in [1]),
        .I4(k5b[41]),
        .I5(\r6/t3/t1/p_0_in [1]),
        .O(\r6/p_0_out [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[41]_i_1__5 
       (.I0(\r7/t0/t2/p_1_in [1]),
        .I1(\r7/t2/t0/p_0_in [1]),
        .I2(\r7/t1/t3/p_1_in [1]),
        .I3(\r7/t1/t3/p_0_in [1]),
        .I4(k6b[41]),
        .I5(\r7/t3/t1/p_0_in [1]),
        .O(\r7/p_0_out [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[41]_i_1__6 
       (.I0(\r8/t0/t2/p_1_in [1]),
        .I1(\r8/t2/t0/p_0_in [1]),
        .I2(\r8/t1/t3/p_1_in [1]),
        .I3(\r8/t1/t3/p_0_in [1]),
        .I4(k7b[41]),
        .I5(\r8/t3/t1/p_0_in [1]),
        .O(\r8/p_0_out [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[41]_i_1__7 
       (.I0(\r9/t0/t2/p_1_in [1]),
        .I1(\r9/t2/t0/p_0_in [1]),
        .I2(\r9/t1/t3/p_1_in [1]),
        .I3(\r9/t1/t3/p_0_in [1]),
        .I4(k8b[41]),
        .I5(\r9/t3/t1/p_0_in [1]),
        .O(\r9/p_0_out [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair365" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[41]_i_1__8 
       (.I0(\a10/k2a [9]),
        .I1(\a10/k4a [9]),
        .I2(\rf/p_1_in [9]),
        .O(\rf/p_4_out [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[42]_i_1 
       (.I0(\r1/t0/t2/p_1_in [2]),
        .I1(\r1/t2/t0/p_0_in [2]),
        .I2(\r1/t1/t3/p_1_in [2]),
        .I3(\r1/t1/t3/p_0_in [2]),
        .I4(k0b[42]),
        .I5(\r1/t3/t1/p_0_in [2]),
        .O(\r1/p_0_out [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[42]_i_1__0 
       (.I0(\r2/t0/t2/p_1_in [2]),
        .I1(\r2/t2/t0/p_0_in [2]),
        .I2(\r2/t1/t3/p_1_in [2]),
        .I3(\r2/t1/t3/p_0_in [2]),
        .I4(k1b[42]),
        .I5(\r2/t3/t1/p_0_in [2]),
        .O(\r2/p_0_out [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[42]_i_1__1 
       (.I0(\r3/t0/t2/p_1_in [2]),
        .I1(\r3/t2/t0/p_0_in [2]),
        .I2(\r3/t1/t3/p_1_in [2]),
        .I3(\r3/t1/t3/p_0_in [2]),
        .I4(k2b[42]),
        .I5(\r3/t3/t1/p_0_in [2]),
        .O(\r3/p_0_out [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[42]_i_1__2 
       (.I0(\r4/t0/t2/p_1_in [2]),
        .I1(\r4/t2/t0/p_0_in [2]),
        .I2(\r4/t1/t3/p_1_in [2]),
        .I3(\r4/t1/t3/p_0_in [2]),
        .I4(k3b[42]),
        .I5(\r4/t3/t1/p_0_in [2]),
        .O(\r4/p_0_out [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[42]_i_1__3 
       (.I0(\r5/t0/t2/p_1_in [2]),
        .I1(\r5/t2/t0/p_0_in [2]),
        .I2(\r5/t1/t3/p_1_in [2]),
        .I3(\r5/t1/t3/p_0_in [2]),
        .I4(k4b[42]),
        .I5(\r5/t3/t1/p_0_in [2]),
        .O(\r5/p_0_out [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[42]_i_1__4 
       (.I0(\r6/t0/t2/p_1_in [2]),
        .I1(\r6/t2/t0/p_0_in [2]),
        .I2(\r6/t1/t3/p_1_in [2]),
        .I3(\r6/t1/t3/p_0_in [2]),
        .I4(k5b[42]),
        .I5(\r6/t3/t1/p_0_in [2]),
        .O(\r6/p_0_out [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[42]_i_1__5 
       (.I0(\r7/t0/t2/p_1_in [2]),
        .I1(\r7/t2/t0/p_0_in [2]),
        .I2(\r7/t1/t3/p_1_in [2]),
        .I3(\r7/t1/t3/p_0_in [2]),
        .I4(k6b[42]),
        .I5(\r7/t3/t1/p_0_in [2]),
        .O(\r7/p_0_out [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[42]_i_1__6 
       (.I0(\r8/t0/t2/p_1_in [2]),
        .I1(\r8/t2/t0/p_0_in [2]),
        .I2(\r8/t1/t3/p_1_in [2]),
        .I3(\r8/t1/t3/p_0_in [2]),
        .I4(k7b[42]),
        .I5(\r8/t3/t1/p_0_in [2]),
        .O(\r8/p_0_out [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[42]_i_1__7 
       (.I0(\r9/t0/t2/p_1_in [2]),
        .I1(\r9/t2/t0/p_0_in [2]),
        .I2(\r9/t1/t3/p_1_in [2]),
        .I3(\r9/t1/t3/p_0_in [2]),
        .I4(k8b[42]),
        .I5(\r9/t3/t1/p_0_in [2]),
        .O(\r9/p_0_out [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair364" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[42]_i_1__8 
       (.I0(\a10/k2a [10]),
        .I1(\a10/k4a [10]),
        .I2(\rf/p_1_in [10]),
        .O(\rf/p_4_out [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[43]_i_1 
       (.I0(\r1/t0/t2/p_1_in [3]),
        .I1(\r1/t2/t0/p_0_in [3]),
        .I2(\r1/t1/t3/p_1_in [3]),
        .I3(\r1/t1/t3/p_0_in [3]),
        .I4(k0b[43]),
        .I5(\r1/t3/t1/p_0_in [3]),
        .O(\r1/p_0_out [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[43]_i_1__0 
       (.I0(\r2/t0/t2/p_1_in [3]),
        .I1(\r2/t2/t0/p_0_in [3]),
        .I2(\r2/t1/t3/p_1_in [3]),
        .I3(\r2/t1/t3/p_0_in [3]),
        .I4(k1b[43]),
        .I5(\r2/t3/t1/p_0_in [3]),
        .O(\r2/p_0_out [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[43]_i_1__1 
       (.I0(\r3/t0/t2/p_1_in [3]),
        .I1(\r3/t2/t0/p_0_in [3]),
        .I2(\r3/t1/t3/p_1_in [3]),
        .I3(\r3/t1/t3/p_0_in [3]),
        .I4(k2b[43]),
        .I5(\r3/t3/t1/p_0_in [3]),
        .O(\r3/p_0_out [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[43]_i_1__2 
       (.I0(\r4/t0/t2/p_1_in [3]),
        .I1(\r4/t2/t0/p_0_in [3]),
        .I2(\r4/t1/t3/p_1_in [3]),
        .I3(\r4/t1/t3/p_0_in [3]),
        .I4(k3b[43]),
        .I5(\r4/t3/t1/p_0_in [3]),
        .O(\r4/p_0_out [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[43]_i_1__3 
       (.I0(\r5/t0/t2/p_1_in [3]),
        .I1(\r5/t2/t0/p_0_in [3]),
        .I2(\r5/t1/t3/p_1_in [3]),
        .I3(\r5/t1/t3/p_0_in [3]),
        .I4(k4b[43]),
        .I5(\r5/t3/t1/p_0_in [3]),
        .O(\r5/p_0_out [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[43]_i_1__4 
       (.I0(\r6/t0/t2/p_1_in [3]),
        .I1(\r6/t2/t0/p_0_in [3]),
        .I2(\r6/t1/t3/p_1_in [3]),
        .I3(\r6/t1/t3/p_0_in [3]),
        .I4(k5b[43]),
        .I5(\r6/t3/t1/p_0_in [3]),
        .O(\r6/p_0_out [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[43]_i_1__5 
       (.I0(\r7/t0/t2/p_1_in [3]),
        .I1(\r7/t2/t0/p_0_in [3]),
        .I2(\r7/t1/t3/p_1_in [3]),
        .I3(\r7/t1/t3/p_0_in [3]),
        .I4(k6b[43]),
        .I5(\r7/t3/t1/p_0_in [3]),
        .O(\r7/p_0_out [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[43]_i_1__6 
       (.I0(\r8/t0/t2/p_1_in [3]),
        .I1(\r8/t2/t0/p_0_in [3]),
        .I2(\r8/t1/t3/p_1_in [3]),
        .I3(\r8/t1/t3/p_0_in [3]),
        .I4(k7b[43]),
        .I5(\r8/t3/t1/p_0_in [3]),
        .O(\r8/p_0_out [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[43]_i_1__7 
       (.I0(\r9/t0/t2/p_1_in [3]),
        .I1(\r9/t2/t0/p_0_in [3]),
        .I2(\r9/t1/t3/p_1_in [3]),
        .I3(\r9/t1/t3/p_0_in [3]),
        .I4(k8b[43]),
        .I5(\r9/t3/t1/p_0_in [3]),
        .O(\r9/p_0_out [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair363" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[43]_i_1__8 
       (.I0(\a10/k2a [11]),
        .I1(\a10/k4a [11]),
        .I2(\rf/p_1_in [11]),
        .O(\rf/p_4_out [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[44]_i_1 
       (.I0(\r1/t0/t2/p_1_in [4]),
        .I1(\r1/t2/t0/p_0_in [4]),
        .I2(\r1/t1/t3/p_1_in [4]),
        .I3(\r1/t1/t3/p_0_in [4]),
        .I4(k0b[44]),
        .I5(\r1/t3/t1/p_0_in [4]),
        .O(\r1/p_0_out [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[44]_i_1__0 
       (.I0(\r2/t0/t2/p_1_in [4]),
        .I1(\r2/t2/t0/p_0_in [4]),
        .I2(\r2/t1/t3/p_1_in [4]),
        .I3(\r2/t1/t3/p_0_in [4]),
        .I4(k1b[44]),
        .I5(\r2/t3/t1/p_0_in [4]),
        .O(\r2/p_0_out [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[44]_i_1__1 
       (.I0(\r3/t0/t2/p_1_in [4]),
        .I1(\r3/t2/t0/p_0_in [4]),
        .I2(\r3/t1/t3/p_1_in [4]),
        .I3(\r3/t1/t3/p_0_in [4]),
        .I4(k2b[44]),
        .I5(\r3/t3/t1/p_0_in [4]),
        .O(\r3/p_0_out [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[44]_i_1__2 
       (.I0(\r4/t0/t2/p_1_in [4]),
        .I1(\r4/t2/t0/p_0_in [4]),
        .I2(\r4/t1/t3/p_1_in [4]),
        .I3(\r4/t1/t3/p_0_in [4]),
        .I4(k3b[44]),
        .I5(\r4/t3/t1/p_0_in [4]),
        .O(\r4/p_0_out [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[44]_i_1__3 
       (.I0(\r5/t0/t2/p_1_in [4]),
        .I1(\r5/t2/t0/p_0_in [4]),
        .I2(\r5/t1/t3/p_1_in [4]),
        .I3(\r5/t1/t3/p_0_in [4]),
        .I4(k4b[44]),
        .I5(\r5/t3/t1/p_0_in [4]),
        .O(\r5/p_0_out [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[44]_i_1__4 
       (.I0(\r6/t0/t2/p_1_in [4]),
        .I1(\r6/t2/t0/p_0_in [4]),
        .I2(\r6/t1/t3/p_1_in [4]),
        .I3(\r6/t1/t3/p_0_in [4]),
        .I4(k5b[44]),
        .I5(\r6/t3/t1/p_0_in [4]),
        .O(\r6/p_0_out [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[44]_i_1__5 
       (.I0(\r7/t0/t2/p_1_in [4]),
        .I1(\r7/t2/t0/p_0_in [4]),
        .I2(\r7/t1/t3/p_1_in [4]),
        .I3(\r7/t1/t3/p_0_in [4]),
        .I4(k6b[44]),
        .I5(\r7/t3/t1/p_0_in [4]),
        .O(\r7/p_0_out [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[44]_i_1__6 
       (.I0(\r8/t0/t2/p_1_in [4]),
        .I1(\r8/t2/t0/p_0_in [4]),
        .I2(\r8/t1/t3/p_1_in [4]),
        .I3(\r8/t1/t3/p_0_in [4]),
        .I4(k7b[44]),
        .I5(\r8/t3/t1/p_0_in [4]),
        .O(\r8/p_0_out [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[44]_i_1__7 
       (.I0(\r9/t0/t2/p_1_in [4]),
        .I1(\r9/t2/t0/p_0_in [4]),
        .I2(\r9/t1/t3/p_1_in [4]),
        .I3(\r9/t1/t3/p_0_in [4]),
        .I4(k8b[44]),
        .I5(\r9/t3/t1/p_0_in [4]),
        .O(\r9/p_0_out [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair362" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[44]_i_1__8 
       (.I0(\a10/k2a [12]),
        .I1(\a10/k4a [12]),
        .I2(\rf/p_1_in [12]),
        .O(\rf/p_4_out [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[45]_i_1 
       (.I0(\r1/t0/t2/p_1_in [5]),
        .I1(\r1/t2/t0/p_0_in [5]),
        .I2(\r1/t1/t3/p_1_in [5]),
        .I3(\r1/t1/t3/p_0_in [5]),
        .I4(k0b[45]),
        .I5(\r1/t3/t1/p_0_in [5]),
        .O(\r1/p_0_out [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[45]_i_1__0 
       (.I0(\r2/t0/t2/p_1_in [5]),
        .I1(\r2/t2/t0/p_0_in [5]),
        .I2(\r2/t1/t3/p_1_in [5]),
        .I3(\r2/t1/t3/p_0_in [5]),
        .I4(k1b[45]),
        .I5(\r2/t3/t1/p_0_in [5]),
        .O(\r2/p_0_out [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[45]_i_1__1 
       (.I0(\r3/t0/t2/p_1_in [5]),
        .I1(\r3/t2/t0/p_0_in [5]),
        .I2(\r3/t1/t3/p_1_in [5]),
        .I3(\r3/t1/t3/p_0_in [5]),
        .I4(k2b[45]),
        .I5(\r3/t3/t1/p_0_in [5]),
        .O(\r3/p_0_out [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[45]_i_1__2 
       (.I0(\r4/t0/t2/p_1_in [5]),
        .I1(\r4/t2/t0/p_0_in [5]),
        .I2(\r4/t1/t3/p_1_in [5]),
        .I3(\r4/t1/t3/p_0_in [5]),
        .I4(k3b[45]),
        .I5(\r4/t3/t1/p_0_in [5]),
        .O(\r4/p_0_out [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[45]_i_1__3 
       (.I0(\r5/t0/t2/p_1_in [5]),
        .I1(\r5/t2/t0/p_0_in [5]),
        .I2(\r5/t1/t3/p_1_in [5]),
        .I3(\r5/t1/t3/p_0_in [5]),
        .I4(k4b[45]),
        .I5(\r5/t3/t1/p_0_in [5]),
        .O(\r5/p_0_out [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[45]_i_1__4 
       (.I0(\r6/t0/t2/p_1_in [5]),
        .I1(\r6/t2/t0/p_0_in [5]),
        .I2(\r6/t1/t3/p_1_in [5]),
        .I3(\r6/t1/t3/p_0_in [5]),
        .I4(k5b[45]),
        .I5(\r6/t3/t1/p_0_in [5]),
        .O(\r6/p_0_out [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[45]_i_1__5 
       (.I0(\r7/t0/t2/p_1_in [5]),
        .I1(\r7/t2/t0/p_0_in [5]),
        .I2(\r7/t1/t3/p_1_in [5]),
        .I3(\r7/t1/t3/p_0_in [5]),
        .I4(k6b[45]),
        .I5(\r7/t3/t1/p_0_in [5]),
        .O(\r7/p_0_out [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[45]_i_1__6 
       (.I0(\r8/t0/t2/p_1_in [5]),
        .I1(\r8/t2/t0/p_0_in [5]),
        .I2(\r8/t1/t3/p_1_in [5]),
        .I3(\r8/t1/t3/p_0_in [5]),
        .I4(k7b[45]),
        .I5(\r8/t3/t1/p_0_in [5]),
        .O(\r8/p_0_out [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[45]_i_1__7 
       (.I0(\r9/t0/t2/p_1_in [5]),
        .I1(\r9/t2/t0/p_0_in [5]),
        .I2(\r9/t1/t3/p_1_in [5]),
        .I3(\r9/t1/t3/p_0_in [5]),
        .I4(k8b[45]),
        .I5(\r9/t3/t1/p_0_in [5]),
        .O(\r9/p_0_out [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair361" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[45]_i_1__8 
       (.I0(\a10/k2a [13]),
        .I1(\a10/k4a [13]),
        .I2(\rf/p_1_in [13]),
        .O(\rf/p_4_out [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[46]_i_1 
       (.I0(\r1/t0/t2/p_1_in [6]),
        .I1(\r1/t2/t0/p_0_in [6]),
        .I2(\r1/t1/t3/p_1_in [6]),
        .I3(\r1/t1/t3/p_0_in [6]),
        .I4(k0b[46]),
        .I5(\r1/t3/t1/p_0_in [6]),
        .O(\r1/p_0_out [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[46]_i_1__0 
       (.I0(\r2/t0/t2/p_1_in [6]),
        .I1(\r2/t2/t0/p_0_in [6]),
        .I2(\r2/t1/t3/p_1_in [6]),
        .I3(\r2/t1/t3/p_0_in [6]),
        .I4(k1b[46]),
        .I5(\r2/t3/t1/p_0_in [6]),
        .O(\r2/p_0_out [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[46]_i_1__1 
       (.I0(\r3/t0/t2/p_1_in [6]),
        .I1(\r3/t2/t0/p_0_in [6]),
        .I2(\r3/t1/t3/p_1_in [6]),
        .I3(\r3/t1/t3/p_0_in [6]),
        .I4(k2b[46]),
        .I5(\r3/t3/t1/p_0_in [6]),
        .O(\r3/p_0_out [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[46]_i_1__2 
       (.I0(\r4/t0/t2/p_1_in [6]),
        .I1(\r4/t2/t0/p_0_in [6]),
        .I2(\r4/t1/t3/p_1_in [6]),
        .I3(\r4/t1/t3/p_0_in [6]),
        .I4(k3b[46]),
        .I5(\r4/t3/t1/p_0_in [6]),
        .O(\r4/p_0_out [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[46]_i_1__3 
       (.I0(\r5/t0/t2/p_1_in [6]),
        .I1(\r5/t2/t0/p_0_in [6]),
        .I2(\r5/t1/t3/p_1_in [6]),
        .I3(\r5/t1/t3/p_0_in [6]),
        .I4(k4b[46]),
        .I5(\r5/t3/t1/p_0_in [6]),
        .O(\r5/p_0_out [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[46]_i_1__4 
       (.I0(\r6/t0/t2/p_1_in [6]),
        .I1(\r6/t2/t0/p_0_in [6]),
        .I2(\r6/t1/t3/p_1_in [6]),
        .I3(\r6/t1/t3/p_0_in [6]),
        .I4(k5b[46]),
        .I5(\r6/t3/t1/p_0_in [6]),
        .O(\r6/p_0_out [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[46]_i_1__5 
       (.I0(\r7/t0/t2/p_1_in [6]),
        .I1(\r7/t2/t0/p_0_in [6]),
        .I2(\r7/t1/t3/p_1_in [6]),
        .I3(\r7/t1/t3/p_0_in [6]),
        .I4(k6b[46]),
        .I5(\r7/t3/t1/p_0_in [6]),
        .O(\r7/p_0_out [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[46]_i_1__6 
       (.I0(\r8/t0/t2/p_1_in [6]),
        .I1(\r8/t2/t0/p_0_in [6]),
        .I2(\r8/t1/t3/p_1_in [6]),
        .I3(\r8/t1/t3/p_0_in [6]),
        .I4(k7b[46]),
        .I5(\r8/t3/t1/p_0_in [6]),
        .O(\r8/p_0_out [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[46]_i_1__7 
       (.I0(\r9/t0/t2/p_1_in [6]),
        .I1(\r9/t2/t0/p_0_in [6]),
        .I2(\r9/t1/t3/p_1_in [6]),
        .I3(\r9/t1/t3/p_0_in [6]),
        .I4(k8b[46]),
        .I5(\r9/t3/t1/p_0_in [6]),
        .O(\r9/p_0_out [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair383" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[46]_i_1__8 
       (.I0(\a10/k2a [14]),
        .I1(\a10/k4a [14]),
        .I2(\rf/p_1_in [14]),
        .O(\rf/p_4_out [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[47]_i_1 
       (.I0(\r1/t0/t2/p_1_in [7]),
        .I1(\r1/t2/t0/p_0_in [7]),
        .I2(\r1/t1/t3/p_1_in [7]),
        .I3(\r1/t1/t3/p_0_in [7]),
        .I4(k0b[47]),
        .I5(\r1/t3/t1/p_0_in [7]),
        .O(\r1/p_0_out [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[47]_i_1__0 
       (.I0(\r2/t0/t2/p_1_in [7]),
        .I1(\r2/t2/t0/p_0_in [7]),
        .I2(\r2/t1/t3/p_1_in [7]),
        .I3(\r2/t1/t3/p_0_in [7]),
        .I4(k1b[47]),
        .I5(\r2/t3/t1/p_0_in [7]),
        .O(\r2/p_0_out [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[47]_i_1__1 
       (.I0(\r3/t0/t2/p_1_in [7]),
        .I1(\r3/t2/t0/p_0_in [7]),
        .I2(\r3/t1/t3/p_1_in [7]),
        .I3(\r3/t1/t3/p_0_in [7]),
        .I4(k2b[47]),
        .I5(\r3/t3/t1/p_0_in [7]),
        .O(\r3/p_0_out [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[47]_i_1__2 
       (.I0(\r4/t0/t2/p_1_in [7]),
        .I1(\r4/t2/t0/p_0_in [7]),
        .I2(\r4/t1/t3/p_1_in [7]),
        .I3(\r4/t1/t3/p_0_in [7]),
        .I4(k3b[47]),
        .I5(\r4/t3/t1/p_0_in [7]),
        .O(\r4/p_0_out [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[47]_i_1__3 
       (.I0(\r5/t0/t2/p_1_in [7]),
        .I1(\r5/t2/t0/p_0_in [7]),
        .I2(\r5/t1/t3/p_1_in [7]),
        .I3(\r5/t1/t3/p_0_in [7]),
        .I4(k4b[47]),
        .I5(\r5/t3/t1/p_0_in [7]),
        .O(\r5/p_0_out [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[47]_i_1__4 
       (.I0(\r6/t0/t2/p_1_in [7]),
        .I1(\r6/t2/t0/p_0_in [7]),
        .I2(\r6/t1/t3/p_1_in [7]),
        .I3(\r6/t1/t3/p_0_in [7]),
        .I4(k5b[47]),
        .I5(\r6/t3/t1/p_0_in [7]),
        .O(\r6/p_0_out [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[47]_i_1__5 
       (.I0(\r7/t0/t2/p_1_in [7]),
        .I1(\r7/t2/t0/p_0_in [7]),
        .I2(\r7/t1/t3/p_1_in [7]),
        .I3(\r7/t1/t3/p_0_in [7]),
        .I4(k6b[47]),
        .I5(\r7/t3/t1/p_0_in [7]),
        .O(\r7/p_0_out [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[47]_i_1__6 
       (.I0(\r8/t0/t2/p_1_in [7]),
        .I1(\r8/t2/t0/p_0_in [7]),
        .I2(\r8/t1/t3/p_1_in [7]),
        .I3(\r8/t1/t3/p_0_in [7]),
        .I4(k7b[47]),
        .I5(\r8/t3/t1/p_0_in [7]),
        .O(\r8/p_0_out [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[47]_i_1__7 
       (.I0(\r9/t0/t2/p_1_in [7]),
        .I1(\r9/t2/t0/p_0_in [7]),
        .I2(\r9/t1/t3/p_1_in [7]),
        .I3(\r9/t1/t3/p_0_in [7]),
        .I4(k8b[47]),
        .I5(\r9/t3/t1/p_0_in [7]),
        .O(\r9/p_0_out [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair382" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[47]_i_1__8 
       (.I0(\a10/k2a [15]),
        .I1(\a10/k4a [15]),
        .I2(\rf/p_1_in [15]),
        .O(\rf/p_4_out [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[48]_i_1 
       (.I0(\r1/t0/t2/p_1_in [0]),
        .I1(\r1/t0/t2/p_0_in [0]),
        .I2(\r1/t2/t0/p_0_in [0]),
        .I3(\r1/t1/t3/p_0_in [0]),
        .I4(k0b[48]),
        .I5(\r1/t3/t1/p_1_in [0]),
        .O(\r1/p_0_out [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[48]_i_1__0 
       (.I0(\r2/t0/t2/p_1_in [0]),
        .I1(\r2/t0/t2/p_0_in [0]),
        .I2(\r2/t2/t0/p_0_in [0]),
        .I3(\r2/t1/t3/p_0_in [0]),
        .I4(k1b[48]),
        .I5(\r2/t3/t1/p_1_in [0]),
        .O(\r2/p_0_out [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[48]_i_1__1 
       (.I0(\r3/t0/t2/p_1_in [0]),
        .I1(\r3/t0/t2/p_0_in [0]),
        .I2(\r3/t2/t0/p_0_in [0]),
        .I3(\r3/t1/t3/p_0_in [0]),
        .I4(k2b[48]),
        .I5(\r3/t3/t1/p_1_in [0]),
        .O(\r3/p_0_out [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[48]_i_1__2 
       (.I0(\r4/t0/t2/p_1_in [0]),
        .I1(\r4/t0/t2/p_0_in [0]),
        .I2(\r4/t2/t0/p_0_in [0]),
        .I3(\r4/t1/t3/p_0_in [0]),
        .I4(k3b[48]),
        .I5(\r4/t3/t1/p_1_in [0]),
        .O(\r4/p_0_out [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[48]_i_1__3 
       (.I0(\r5/t0/t2/p_1_in [0]),
        .I1(\r5/t0/t2/p_0_in [0]),
        .I2(\r5/t2/t0/p_0_in [0]),
        .I3(\r5/t1/t3/p_0_in [0]),
        .I4(k4b[48]),
        .I5(\r5/t3/t1/p_1_in [0]),
        .O(\r5/p_0_out [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[48]_i_1__4 
       (.I0(\r6/t0/t2/p_1_in [0]),
        .I1(\r6/t0/t2/p_0_in [0]),
        .I2(\r6/t2/t0/p_0_in [0]),
        .I3(\r6/t1/t3/p_0_in [0]),
        .I4(k5b[48]),
        .I5(\r6/t3/t1/p_1_in [0]),
        .O(\r6/p_0_out [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[48]_i_1__5 
       (.I0(\r7/t0/t2/p_1_in [0]),
        .I1(\r7/t0/t2/p_0_in [0]),
        .I2(\r7/t2/t0/p_0_in [0]),
        .I3(\r7/t1/t3/p_0_in [0]),
        .I4(k6b[48]),
        .I5(\r7/t3/t1/p_1_in [0]),
        .O(\r7/p_0_out [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[48]_i_1__6 
       (.I0(\r8/t0/t2/p_1_in [0]),
        .I1(\r8/t0/t2/p_0_in [0]),
        .I2(\r8/t2/t0/p_0_in [0]),
        .I3(\r8/t1/t3/p_0_in [0]),
        .I4(k7b[48]),
        .I5(\r8/t3/t1/p_1_in [0]),
        .O(\r8/p_0_out [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[48]_i_1__7 
       (.I0(\r9/t0/t2/p_1_in [0]),
        .I1(\r9/t0/t2/p_0_in [0]),
        .I2(\r9/t2/t0/p_0_in [0]),
        .I3(\r9/t1/t3/p_0_in [0]),
        .I4(k8b[48]),
        .I5(\r9/t3/t1/p_1_in [0]),
        .O(\r9/p_0_out [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair381" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[48]_i_1__8 
       (.I0(\a10/k2a [16]),
        .I1(\a10/k4a [16]),
        .I2(\rf/p_1_in [16]),
        .O(\rf/p_4_out [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[49]_i_1 
       (.I0(\r1/t0/t2/p_1_in [1]),
        .I1(\r1/t0/t2/p_0_in [1]),
        .I2(\r1/t2/t0/p_0_in [1]),
        .I3(\r1/t1/t3/p_0_in [1]),
        .I4(k0b[49]),
        .I5(\r1/t3/t1/p_1_in [1]),
        .O(\r1/p_0_out [49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[49]_i_1__0 
       (.I0(\r2/t0/t2/p_1_in [1]),
        .I1(\r2/t0/t2/p_0_in [1]),
        .I2(\r2/t2/t0/p_0_in [1]),
        .I3(\r2/t1/t3/p_0_in [1]),
        .I4(k1b[49]),
        .I5(\r2/t3/t1/p_1_in [1]),
        .O(\r2/p_0_out [49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[49]_i_1__1 
       (.I0(\r3/t0/t2/p_1_in [1]),
        .I1(\r3/t0/t2/p_0_in [1]),
        .I2(\r3/t2/t0/p_0_in [1]),
        .I3(\r3/t1/t3/p_0_in [1]),
        .I4(k2b[49]),
        .I5(\r3/t3/t1/p_1_in [1]),
        .O(\r3/p_0_out [49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[49]_i_1__2 
       (.I0(\r4/t0/t2/p_1_in [1]),
        .I1(\r4/t0/t2/p_0_in [1]),
        .I2(\r4/t2/t0/p_0_in [1]),
        .I3(\r4/t1/t3/p_0_in [1]),
        .I4(k3b[49]),
        .I5(\r4/t3/t1/p_1_in [1]),
        .O(\r4/p_0_out [49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[49]_i_1__3 
       (.I0(\r5/t0/t2/p_1_in [1]),
        .I1(\r5/t0/t2/p_0_in [1]),
        .I2(\r5/t2/t0/p_0_in [1]),
        .I3(\r5/t1/t3/p_0_in [1]),
        .I4(k4b[49]),
        .I5(\r5/t3/t1/p_1_in [1]),
        .O(\r5/p_0_out [49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[49]_i_1__4 
       (.I0(\r6/t0/t2/p_1_in [1]),
        .I1(\r6/t0/t2/p_0_in [1]),
        .I2(\r6/t2/t0/p_0_in [1]),
        .I3(\r6/t1/t3/p_0_in [1]),
        .I4(k5b[49]),
        .I5(\r6/t3/t1/p_1_in [1]),
        .O(\r6/p_0_out [49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[49]_i_1__5 
       (.I0(\r7/t0/t2/p_1_in [1]),
        .I1(\r7/t0/t2/p_0_in [1]),
        .I2(\r7/t2/t0/p_0_in [1]),
        .I3(\r7/t1/t3/p_0_in [1]),
        .I4(k6b[49]),
        .I5(\r7/t3/t1/p_1_in [1]),
        .O(\r7/p_0_out [49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[49]_i_1__6 
       (.I0(\r8/t0/t2/p_1_in [1]),
        .I1(\r8/t0/t2/p_0_in [1]),
        .I2(\r8/t2/t0/p_0_in [1]),
        .I3(\r8/t1/t3/p_0_in [1]),
        .I4(k7b[49]),
        .I5(\r8/t3/t1/p_1_in [1]),
        .O(\r8/p_0_out [49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[49]_i_1__7 
       (.I0(\r9/t0/t2/p_1_in [1]),
        .I1(\r9/t0/t2/p_0_in [1]),
        .I2(\r9/t2/t0/p_0_in [1]),
        .I3(\r9/t1/t3/p_0_in [1]),
        .I4(k8b[49]),
        .I5(\r9/t3/t1/p_1_in [1]),
        .O(\r9/p_0_out [49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair380" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[49]_i_1__8 
       (.I0(\a10/k2a [17]),
        .I1(\a10/k4a [17]),
        .I2(\rf/p_1_in [17]),
        .O(\rf/p_4_out [49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[4]_i_1 
       (.I0(\r1/t0/t1/p_0_in [4]),
        .I1(\r1/t2/t3/p_1_in [4]),
        .I2(\r1/t1/t2/p_0_in [4]),
        .I3(k0b[4]),
        .I4(\r1/t3/t0/p_1_in [4]),
        .I5(\r1/t3/t0/p_0_in [4]),
        .O(\r1/p_0_out [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[4]_i_1__0 
       (.I0(\r2/t0/t1/p_0_in [4]),
        .I1(\r2/t2/t3/p_1_in [4]),
        .I2(\r2/t1/t2/p_0_in [4]),
        .I3(k1b[4]),
        .I4(\r2/t3/t0/p_1_in [4]),
        .I5(\r2/t3/t0/p_0_in [4]),
        .O(\r2/p_0_out [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[4]_i_1__1 
       (.I0(\r3/t0/t1/p_0_in [4]),
        .I1(\r3/t2/t3/p_1_in [4]),
        .I2(\r3/t1/t2/p_0_in [4]),
        .I3(k2b[4]),
        .I4(\r3/t3/t0/p_1_in [4]),
        .I5(\r3/t3/t0/p_0_in [4]),
        .O(\r3/p_0_out [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[4]_i_1__2 
       (.I0(\r4/t0/t1/p_0_in [4]),
        .I1(\r4/t2/t3/p_1_in [4]),
        .I2(\r4/t1/t2/p_0_in [4]),
        .I3(k3b[4]),
        .I4(\r4/t3/t0/p_1_in [4]),
        .I5(\r4/t3/t0/p_0_in [4]),
        .O(\r4/p_0_out [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[4]_i_1__3 
       (.I0(\r5/t0/t1/p_0_in [4]),
        .I1(\r5/t2/t3/p_1_in [4]),
        .I2(\r5/t1/t2/p_0_in [4]),
        .I3(k4b[4]),
        .I4(\r5/t3/t0/p_1_in [4]),
        .I5(\r5/t3/t0/p_0_in [4]),
        .O(\r5/p_0_out [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[4]_i_1__4 
       (.I0(\r6/t0/t1/p_0_in [4]),
        .I1(\r6/t2/t3/p_1_in [4]),
        .I2(\r6/t1/t2/p_0_in [4]),
        .I3(k5b[4]),
        .I4(\r6/t3/t0/p_1_in [4]),
        .I5(\r6/t3/t0/p_0_in [4]),
        .O(\r6/p_0_out [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[4]_i_1__5 
       (.I0(\r7/t0/t1/p_0_in [4]),
        .I1(\r7/t2/t3/p_1_in [4]),
        .I2(\r7/t1/t2/p_0_in [4]),
        .I3(k6b[4]),
        .I4(\r7/t3/t0/p_1_in [4]),
        .I5(\r7/t3/t0/p_0_in [4]),
        .O(\r7/p_0_out [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[4]_i_1__6 
       (.I0(\r8/t0/t1/p_0_in [4]),
        .I1(\r8/t2/t3/p_1_in [4]),
        .I2(\r8/t1/t2/p_0_in [4]),
        .I3(k7b[4]),
        .I4(\r8/t3/t0/p_1_in [4]),
        .I5(\r8/t3/t0/p_0_in [4]),
        .O(\r8/p_0_out [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[4]_i_1__7 
       (.I0(\r9/t0/t1/p_0_in [4]),
        .I1(\r9/t2/t3/p_1_in [4]),
        .I2(\r9/t1/t2/p_0_in [4]),
        .I3(k8b[4]),
        .I4(\r9/t3/t0/p_1_in [4]),
        .I5(\r9/t3/t0/p_0_in [4]),
        .O(\r9/p_0_out [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair338" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[4]_i_1__8 
       (.I0(\a10/k3a [4]),
        .I1(\a10/k4a [4]),
        .I2(\rf/p_0_in [4]),
        .O(\rf/p_4_out [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[50]_i_1 
       (.I0(\r1/t0/t2/p_1_in [2]),
        .I1(\r1/t0/t2/p_0_in [2]),
        .I2(\r1/t2/t0/p_0_in [2]),
        .I3(\r1/t1/t3/p_0_in [2]),
        .I4(k0b[50]),
        .I5(\r1/t3/t1/p_1_in [2]),
        .O(\r1/p_0_out [50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[50]_i_1__0 
       (.I0(\r2/t0/t2/p_1_in [2]),
        .I1(\r2/t0/t2/p_0_in [2]),
        .I2(\r2/t2/t0/p_0_in [2]),
        .I3(\r2/t1/t3/p_0_in [2]),
        .I4(k1b[50]),
        .I5(\r2/t3/t1/p_1_in [2]),
        .O(\r2/p_0_out [50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[50]_i_1__1 
       (.I0(\r3/t0/t2/p_1_in [2]),
        .I1(\r3/t0/t2/p_0_in [2]),
        .I2(\r3/t2/t0/p_0_in [2]),
        .I3(\r3/t1/t3/p_0_in [2]),
        .I4(k2b[50]),
        .I5(\r3/t3/t1/p_1_in [2]),
        .O(\r3/p_0_out [50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[50]_i_1__2 
       (.I0(\r4/t0/t2/p_1_in [2]),
        .I1(\r4/t0/t2/p_0_in [2]),
        .I2(\r4/t2/t0/p_0_in [2]),
        .I3(\r4/t1/t3/p_0_in [2]),
        .I4(k3b[50]),
        .I5(\r4/t3/t1/p_1_in [2]),
        .O(\r4/p_0_out [50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[50]_i_1__3 
       (.I0(\r5/t0/t2/p_1_in [2]),
        .I1(\r5/t0/t2/p_0_in [2]),
        .I2(\r5/t2/t0/p_0_in [2]),
        .I3(\r5/t1/t3/p_0_in [2]),
        .I4(k4b[50]),
        .I5(\r5/t3/t1/p_1_in [2]),
        .O(\r5/p_0_out [50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[50]_i_1__4 
       (.I0(\r6/t0/t2/p_1_in [2]),
        .I1(\r6/t0/t2/p_0_in [2]),
        .I2(\r6/t2/t0/p_0_in [2]),
        .I3(\r6/t1/t3/p_0_in [2]),
        .I4(k5b[50]),
        .I5(\r6/t3/t1/p_1_in [2]),
        .O(\r6/p_0_out [50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[50]_i_1__5 
       (.I0(\r7/t0/t2/p_1_in [2]),
        .I1(\r7/t0/t2/p_0_in [2]),
        .I2(\r7/t2/t0/p_0_in [2]),
        .I3(\r7/t1/t3/p_0_in [2]),
        .I4(k6b[50]),
        .I5(\r7/t3/t1/p_1_in [2]),
        .O(\r7/p_0_out [50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[50]_i_1__6 
       (.I0(\r8/t0/t2/p_1_in [2]),
        .I1(\r8/t0/t2/p_0_in [2]),
        .I2(\r8/t2/t0/p_0_in [2]),
        .I3(\r8/t1/t3/p_0_in [2]),
        .I4(k7b[50]),
        .I5(\r8/t3/t1/p_1_in [2]),
        .O(\r8/p_0_out [50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[50]_i_1__7 
       (.I0(\r9/t0/t2/p_1_in [2]),
        .I1(\r9/t0/t2/p_0_in [2]),
        .I2(\r9/t2/t0/p_0_in [2]),
        .I3(\r9/t1/t3/p_0_in [2]),
        .I4(k8b[50]),
        .I5(\r9/t3/t1/p_1_in [2]),
        .O(\r9/p_0_out [50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair379" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[50]_i_1__8 
       (.I0(\a10/k2a [18]),
        .I1(\a10/k4a [18]),
        .I2(\rf/p_1_in [18]),
        .O(\rf/p_4_out [50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[51]_i_1 
       (.I0(\r1/t0/t2/p_1_in [3]),
        .I1(\r1/t0/t2/p_0_in [3]),
        .I2(\r1/t2/t0/p_0_in [3]),
        .I3(\r1/t1/t3/p_0_in [3]),
        .I4(k0b[51]),
        .I5(\r1/t3/t1/p_1_in [3]),
        .O(\r1/p_0_out [51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[51]_i_1__0 
       (.I0(\r2/t0/t2/p_1_in [3]),
        .I1(\r2/t0/t2/p_0_in [3]),
        .I2(\r2/t2/t0/p_0_in [3]),
        .I3(\r2/t1/t3/p_0_in [3]),
        .I4(k1b[51]),
        .I5(\r2/t3/t1/p_1_in [3]),
        .O(\r2/p_0_out [51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[51]_i_1__1 
       (.I0(\r3/t0/t2/p_1_in [3]),
        .I1(\r3/t0/t2/p_0_in [3]),
        .I2(\r3/t2/t0/p_0_in [3]),
        .I3(\r3/t1/t3/p_0_in [3]),
        .I4(k2b[51]),
        .I5(\r3/t3/t1/p_1_in [3]),
        .O(\r3/p_0_out [51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[51]_i_1__2 
       (.I0(\r4/t0/t2/p_1_in [3]),
        .I1(\r4/t0/t2/p_0_in [3]),
        .I2(\r4/t2/t0/p_0_in [3]),
        .I3(\r4/t1/t3/p_0_in [3]),
        .I4(k3b[51]),
        .I5(\r4/t3/t1/p_1_in [3]),
        .O(\r4/p_0_out [51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[51]_i_1__3 
       (.I0(\r5/t0/t2/p_1_in [3]),
        .I1(\r5/t0/t2/p_0_in [3]),
        .I2(\r5/t2/t0/p_0_in [3]),
        .I3(\r5/t1/t3/p_0_in [3]),
        .I4(k4b[51]),
        .I5(\r5/t3/t1/p_1_in [3]),
        .O(\r5/p_0_out [51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[51]_i_1__4 
       (.I0(\r6/t0/t2/p_1_in [3]),
        .I1(\r6/t0/t2/p_0_in [3]),
        .I2(\r6/t2/t0/p_0_in [3]),
        .I3(\r6/t1/t3/p_0_in [3]),
        .I4(k5b[51]),
        .I5(\r6/t3/t1/p_1_in [3]),
        .O(\r6/p_0_out [51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[51]_i_1__5 
       (.I0(\r7/t0/t2/p_1_in [3]),
        .I1(\r7/t0/t2/p_0_in [3]),
        .I2(\r7/t2/t0/p_0_in [3]),
        .I3(\r7/t1/t3/p_0_in [3]),
        .I4(k6b[51]),
        .I5(\r7/t3/t1/p_1_in [3]),
        .O(\r7/p_0_out [51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[51]_i_1__6 
       (.I0(\r8/t0/t2/p_1_in [3]),
        .I1(\r8/t0/t2/p_0_in [3]),
        .I2(\r8/t2/t0/p_0_in [3]),
        .I3(\r8/t1/t3/p_0_in [3]),
        .I4(k7b[51]),
        .I5(\r8/t3/t1/p_1_in [3]),
        .O(\r8/p_0_out [51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[51]_i_1__7 
       (.I0(\r9/t0/t2/p_1_in [3]),
        .I1(\r9/t0/t2/p_0_in [3]),
        .I2(\r9/t2/t0/p_0_in [3]),
        .I3(\r9/t1/t3/p_0_in [3]),
        .I4(k8b[51]),
        .I5(\r9/t3/t1/p_1_in [3]),
        .O(\r9/p_0_out [51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair378" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[51]_i_1__8 
       (.I0(\a10/k2a [19]),
        .I1(\a10/k4a [19]),
        .I2(\rf/p_1_in [19]),
        .O(\rf/p_4_out [51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[52]_i_1 
       (.I0(\r1/t0/t2/p_1_in [4]),
        .I1(\r1/t0/t2/p_0_in [4]),
        .I2(\r1/t2/t0/p_0_in [4]),
        .I3(\r1/t1/t3/p_0_in [4]),
        .I4(k0b[52]),
        .I5(\r1/t3/t1/p_1_in [4]),
        .O(\r1/p_0_out [52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[52]_i_1__0 
       (.I0(\r2/t0/t2/p_1_in [4]),
        .I1(\r2/t0/t2/p_0_in [4]),
        .I2(\r2/t2/t0/p_0_in [4]),
        .I3(\r2/t1/t3/p_0_in [4]),
        .I4(k1b[52]),
        .I5(\r2/t3/t1/p_1_in [4]),
        .O(\r2/p_0_out [52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[52]_i_1__1 
       (.I0(\r3/t0/t2/p_1_in [4]),
        .I1(\r3/t0/t2/p_0_in [4]),
        .I2(\r3/t2/t0/p_0_in [4]),
        .I3(\r3/t1/t3/p_0_in [4]),
        .I4(k2b[52]),
        .I5(\r3/t3/t1/p_1_in [4]),
        .O(\r3/p_0_out [52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[52]_i_1__2 
       (.I0(\r4/t0/t2/p_1_in [4]),
        .I1(\r4/t0/t2/p_0_in [4]),
        .I2(\r4/t2/t0/p_0_in [4]),
        .I3(\r4/t1/t3/p_0_in [4]),
        .I4(k3b[52]),
        .I5(\r4/t3/t1/p_1_in [4]),
        .O(\r4/p_0_out [52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[52]_i_1__3 
       (.I0(\r5/t0/t2/p_1_in [4]),
        .I1(\r5/t0/t2/p_0_in [4]),
        .I2(\r5/t2/t0/p_0_in [4]),
        .I3(\r5/t1/t3/p_0_in [4]),
        .I4(k4b[52]),
        .I5(\r5/t3/t1/p_1_in [4]),
        .O(\r5/p_0_out [52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[52]_i_1__4 
       (.I0(\r6/t0/t2/p_1_in [4]),
        .I1(\r6/t0/t2/p_0_in [4]),
        .I2(\r6/t2/t0/p_0_in [4]),
        .I3(\r6/t1/t3/p_0_in [4]),
        .I4(k5b[52]),
        .I5(\r6/t3/t1/p_1_in [4]),
        .O(\r6/p_0_out [52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[52]_i_1__5 
       (.I0(\r7/t0/t2/p_1_in [4]),
        .I1(\r7/t0/t2/p_0_in [4]),
        .I2(\r7/t2/t0/p_0_in [4]),
        .I3(\r7/t1/t3/p_0_in [4]),
        .I4(k6b[52]),
        .I5(\r7/t3/t1/p_1_in [4]),
        .O(\r7/p_0_out [52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[52]_i_1__6 
       (.I0(\r8/t0/t2/p_1_in [4]),
        .I1(\r8/t0/t2/p_0_in [4]),
        .I2(\r8/t2/t0/p_0_in [4]),
        .I3(\r8/t1/t3/p_0_in [4]),
        .I4(k7b[52]),
        .I5(\r8/t3/t1/p_1_in [4]),
        .O(\r8/p_0_out [52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[52]_i_1__7 
       (.I0(\r9/t0/t2/p_1_in [4]),
        .I1(\r9/t0/t2/p_0_in [4]),
        .I2(\r9/t2/t0/p_0_in [4]),
        .I3(\r9/t1/t3/p_0_in [4]),
        .I4(k8b[52]),
        .I5(\r9/t3/t1/p_1_in [4]),
        .O(\r9/p_0_out [52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair377" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[52]_i_1__8 
       (.I0(\a10/k2a [20]),
        .I1(\a10/k4a [20]),
        .I2(\rf/p_1_in [20]),
        .O(\rf/p_4_out [52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[53]_i_1 
       (.I0(\r1/t0/t2/p_1_in [5]),
        .I1(\r1/t0/t2/p_0_in [5]),
        .I2(\r1/t2/t0/p_0_in [5]),
        .I3(\r1/t1/t3/p_0_in [5]),
        .I4(k0b[53]),
        .I5(\r1/t3/t1/p_1_in [5]),
        .O(\r1/p_0_out [53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[53]_i_1__0 
       (.I0(\r2/t0/t2/p_1_in [5]),
        .I1(\r2/t0/t2/p_0_in [5]),
        .I2(\r2/t2/t0/p_0_in [5]),
        .I3(\r2/t1/t3/p_0_in [5]),
        .I4(k1b[53]),
        .I5(\r2/t3/t1/p_1_in [5]),
        .O(\r2/p_0_out [53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[53]_i_1__1 
       (.I0(\r3/t0/t2/p_1_in [5]),
        .I1(\r3/t0/t2/p_0_in [5]),
        .I2(\r3/t2/t0/p_0_in [5]),
        .I3(\r3/t1/t3/p_0_in [5]),
        .I4(k2b[53]),
        .I5(\r3/t3/t1/p_1_in [5]),
        .O(\r3/p_0_out [53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[53]_i_1__2 
       (.I0(\r4/t0/t2/p_1_in [5]),
        .I1(\r4/t0/t2/p_0_in [5]),
        .I2(\r4/t2/t0/p_0_in [5]),
        .I3(\r4/t1/t3/p_0_in [5]),
        .I4(k3b[53]),
        .I5(\r4/t3/t1/p_1_in [5]),
        .O(\r4/p_0_out [53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[53]_i_1__3 
       (.I0(\r5/t0/t2/p_1_in [5]),
        .I1(\r5/t0/t2/p_0_in [5]),
        .I2(\r5/t2/t0/p_0_in [5]),
        .I3(\r5/t1/t3/p_0_in [5]),
        .I4(k4b[53]),
        .I5(\r5/t3/t1/p_1_in [5]),
        .O(\r5/p_0_out [53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[53]_i_1__4 
       (.I0(\r6/t0/t2/p_1_in [5]),
        .I1(\r6/t0/t2/p_0_in [5]),
        .I2(\r6/t2/t0/p_0_in [5]),
        .I3(\r6/t1/t3/p_0_in [5]),
        .I4(k5b[53]),
        .I5(\r6/t3/t1/p_1_in [5]),
        .O(\r6/p_0_out [53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[53]_i_1__5 
       (.I0(\r7/t0/t2/p_1_in [5]),
        .I1(\r7/t0/t2/p_0_in [5]),
        .I2(\r7/t2/t0/p_0_in [5]),
        .I3(\r7/t1/t3/p_0_in [5]),
        .I4(k6b[53]),
        .I5(\r7/t3/t1/p_1_in [5]),
        .O(\r7/p_0_out [53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[53]_i_1__6 
       (.I0(\r8/t0/t2/p_1_in [5]),
        .I1(\r8/t0/t2/p_0_in [5]),
        .I2(\r8/t2/t0/p_0_in [5]),
        .I3(\r8/t1/t3/p_0_in [5]),
        .I4(k7b[53]),
        .I5(\r8/t3/t1/p_1_in [5]),
        .O(\r8/p_0_out [53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[53]_i_1__7 
       (.I0(\r9/t0/t2/p_1_in [5]),
        .I1(\r9/t0/t2/p_0_in [5]),
        .I2(\r9/t2/t0/p_0_in [5]),
        .I3(\r9/t1/t3/p_0_in [5]),
        .I4(k8b[53]),
        .I5(\r9/t3/t1/p_1_in [5]),
        .O(\r9/p_0_out [53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair376" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[53]_i_1__8 
       (.I0(\a10/k2a [21]),
        .I1(\a10/k4a [21]),
        .I2(\rf/p_1_in [21]),
        .O(\rf/p_4_out [53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[54]_i_1 
       (.I0(\r1/t0/t2/p_1_in [6]),
        .I1(\r1/t0/t2/p_0_in [6]),
        .I2(\r1/t2/t0/p_0_in [6]),
        .I3(\r1/t1/t3/p_0_in [6]),
        .I4(k0b[54]),
        .I5(\r1/t3/t1/p_1_in [6]),
        .O(\r1/p_0_out [54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[54]_i_1__0 
       (.I0(\r2/t0/t2/p_1_in [6]),
        .I1(\r2/t0/t2/p_0_in [6]),
        .I2(\r2/t2/t0/p_0_in [6]),
        .I3(\r2/t1/t3/p_0_in [6]),
        .I4(k1b[54]),
        .I5(\r2/t3/t1/p_1_in [6]),
        .O(\r2/p_0_out [54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[54]_i_1__1 
       (.I0(\r3/t0/t2/p_1_in [6]),
        .I1(\r3/t0/t2/p_0_in [6]),
        .I2(\r3/t2/t0/p_0_in [6]),
        .I3(\r3/t1/t3/p_0_in [6]),
        .I4(k2b[54]),
        .I5(\r3/t3/t1/p_1_in [6]),
        .O(\r3/p_0_out [54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[54]_i_1__2 
       (.I0(\r4/t0/t2/p_1_in [6]),
        .I1(\r4/t0/t2/p_0_in [6]),
        .I2(\r4/t2/t0/p_0_in [6]),
        .I3(\r4/t1/t3/p_0_in [6]),
        .I4(k3b[54]),
        .I5(\r4/t3/t1/p_1_in [6]),
        .O(\r4/p_0_out [54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[54]_i_1__3 
       (.I0(\r5/t0/t2/p_1_in [6]),
        .I1(\r5/t0/t2/p_0_in [6]),
        .I2(\r5/t2/t0/p_0_in [6]),
        .I3(\r5/t1/t3/p_0_in [6]),
        .I4(k4b[54]),
        .I5(\r5/t3/t1/p_1_in [6]),
        .O(\r5/p_0_out [54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[54]_i_1__4 
       (.I0(\r6/t0/t2/p_1_in [6]),
        .I1(\r6/t0/t2/p_0_in [6]),
        .I2(\r6/t2/t0/p_0_in [6]),
        .I3(\r6/t1/t3/p_0_in [6]),
        .I4(k5b[54]),
        .I5(\r6/t3/t1/p_1_in [6]),
        .O(\r6/p_0_out [54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[54]_i_1__5 
       (.I0(\r7/t0/t2/p_1_in [6]),
        .I1(\r7/t0/t2/p_0_in [6]),
        .I2(\r7/t2/t0/p_0_in [6]),
        .I3(\r7/t1/t3/p_0_in [6]),
        .I4(k6b[54]),
        .I5(\r7/t3/t1/p_1_in [6]),
        .O(\r7/p_0_out [54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[54]_i_1__6 
       (.I0(\r8/t0/t2/p_1_in [6]),
        .I1(\r8/t0/t2/p_0_in [6]),
        .I2(\r8/t2/t0/p_0_in [6]),
        .I3(\r8/t1/t3/p_0_in [6]),
        .I4(k7b[54]),
        .I5(\r8/t3/t1/p_1_in [6]),
        .O(\r8/p_0_out [54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[54]_i_1__7 
       (.I0(\r9/t0/t2/p_1_in [6]),
        .I1(\r9/t0/t2/p_0_in [6]),
        .I2(\r9/t2/t0/p_0_in [6]),
        .I3(\r9/t1/t3/p_0_in [6]),
        .I4(k8b[54]),
        .I5(\r9/t3/t1/p_1_in [6]),
        .O(\r9/p_0_out [54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair375" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[54]_i_1__8 
       (.I0(\a10/k2a [22]),
        .I1(\a10/k4a [22]),
        .I2(\rf/p_1_in [22]),
        .O(\rf/p_4_out [54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[55]_i_1 
       (.I0(\r1/t0/t2/p_1_in [7]),
        .I1(\r1/t0/t2/p_0_in [7]),
        .I2(\r1/t2/t0/p_0_in [7]),
        .I3(\r1/t1/t3/p_0_in [7]),
        .I4(k0b[55]),
        .I5(\r1/t3/t1/p_1_in [7]),
        .O(\r1/p_0_out [55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[55]_i_1__0 
       (.I0(\r2/t0/t2/p_1_in [7]),
        .I1(\r2/t0/t2/p_0_in [7]),
        .I2(\r2/t2/t0/p_0_in [7]),
        .I3(\r2/t1/t3/p_0_in [7]),
        .I4(k1b[55]),
        .I5(\r2/t3/t1/p_1_in [7]),
        .O(\r2/p_0_out [55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[55]_i_1__1 
       (.I0(\r3/t0/t2/p_1_in [7]),
        .I1(\r3/t0/t2/p_0_in [7]),
        .I2(\r3/t2/t0/p_0_in [7]),
        .I3(\r3/t1/t3/p_0_in [7]),
        .I4(k2b[55]),
        .I5(\r3/t3/t1/p_1_in [7]),
        .O(\r3/p_0_out [55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[55]_i_1__2 
       (.I0(\r4/t0/t2/p_1_in [7]),
        .I1(\r4/t0/t2/p_0_in [7]),
        .I2(\r4/t2/t0/p_0_in [7]),
        .I3(\r4/t1/t3/p_0_in [7]),
        .I4(k3b[55]),
        .I5(\r4/t3/t1/p_1_in [7]),
        .O(\r4/p_0_out [55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[55]_i_1__3 
       (.I0(\r5/t0/t2/p_1_in [7]),
        .I1(\r5/t0/t2/p_0_in [7]),
        .I2(\r5/t2/t0/p_0_in [7]),
        .I3(\r5/t1/t3/p_0_in [7]),
        .I4(k4b[55]),
        .I5(\r5/t3/t1/p_1_in [7]),
        .O(\r5/p_0_out [55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[55]_i_1__4 
       (.I0(\r6/t0/t2/p_1_in [7]),
        .I1(\r6/t0/t2/p_0_in [7]),
        .I2(\r6/t2/t0/p_0_in [7]),
        .I3(\r6/t1/t3/p_0_in [7]),
        .I4(k5b[55]),
        .I5(\r6/t3/t1/p_1_in [7]),
        .O(\r6/p_0_out [55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[55]_i_1__5 
       (.I0(\r7/t0/t2/p_1_in [7]),
        .I1(\r7/t0/t2/p_0_in [7]),
        .I2(\r7/t2/t0/p_0_in [7]),
        .I3(\r7/t1/t3/p_0_in [7]),
        .I4(k6b[55]),
        .I5(\r7/t3/t1/p_1_in [7]),
        .O(\r7/p_0_out [55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[55]_i_1__6 
       (.I0(\r8/t0/t2/p_1_in [7]),
        .I1(\r8/t0/t2/p_0_in [7]),
        .I2(\r8/t2/t0/p_0_in [7]),
        .I3(\r8/t1/t3/p_0_in [7]),
        .I4(k7b[55]),
        .I5(\r8/t3/t1/p_1_in [7]),
        .O(\r8/p_0_out [55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[55]_i_1__7 
       (.I0(\r9/t0/t2/p_1_in [7]),
        .I1(\r9/t0/t2/p_0_in [7]),
        .I2(\r9/t2/t0/p_0_in [7]),
        .I3(\r9/t1/t3/p_0_in [7]),
        .I4(k8b[55]),
        .I5(\r9/t3/t1/p_1_in [7]),
        .O(\r9/p_0_out [55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair360" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[55]_i_1__8 
       (.I0(\a10/k2a [23]),
        .I1(\a10/k4a [23]),
        .I2(\rf/p_1_in [23]),
        .O(\rf/p_4_out [55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[56]_i_1 
       (.I0(\r1/t0/t2/p_0_in [0]),
        .I1(\r1/t2/t0/p_1_in [0]),
        .I2(\r1/t1/t3/p_0_in [0]),
        .I3(k0b[56]),
        .I4(\r1/t3/t1/p_1_in [0]),
        .I5(\r1/t3/t1/p_0_in [0]),
        .O(\r1/p_0_out [56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[56]_i_1__0 
       (.I0(\r2/t0/t2/p_0_in [0]),
        .I1(\r2/t2/t0/p_1_in [0]),
        .I2(\r2/t1/t3/p_0_in [0]),
        .I3(k1b[56]),
        .I4(\r2/t3/t1/p_1_in [0]),
        .I5(\r2/t3/t1/p_0_in [0]),
        .O(\r2/p_0_out [56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[56]_i_1__1 
       (.I0(\r3/t0/t2/p_0_in [0]),
        .I1(\r3/t2/t0/p_1_in [0]),
        .I2(\r3/t1/t3/p_0_in [0]),
        .I3(k2b[56]),
        .I4(\r3/t3/t1/p_1_in [0]),
        .I5(\r3/t3/t1/p_0_in [0]),
        .O(\r3/p_0_out [56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[56]_i_1__2 
       (.I0(\r4/t0/t2/p_0_in [0]),
        .I1(\r4/t2/t0/p_1_in [0]),
        .I2(\r4/t1/t3/p_0_in [0]),
        .I3(k3b[56]),
        .I4(\r4/t3/t1/p_1_in [0]),
        .I5(\r4/t3/t1/p_0_in [0]),
        .O(\r4/p_0_out [56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[56]_i_1__3 
       (.I0(\r5/t0/t2/p_0_in [0]),
        .I1(\r5/t2/t0/p_1_in [0]),
        .I2(\r5/t1/t3/p_0_in [0]),
        .I3(k4b[56]),
        .I4(\r5/t3/t1/p_1_in [0]),
        .I5(\r5/t3/t1/p_0_in [0]),
        .O(\r5/p_0_out [56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[56]_i_1__4 
       (.I0(\r6/t0/t2/p_0_in [0]),
        .I1(\r6/t2/t0/p_1_in [0]),
        .I2(\r6/t1/t3/p_0_in [0]),
        .I3(k5b[56]),
        .I4(\r6/t3/t1/p_1_in [0]),
        .I5(\r6/t3/t1/p_0_in [0]),
        .O(\r6/p_0_out [56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[56]_i_1__5 
       (.I0(\r7/t0/t2/p_0_in [0]),
        .I1(\r7/t2/t0/p_1_in [0]),
        .I2(\r7/t1/t3/p_0_in [0]),
        .I3(k6b[56]),
        .I4(\r7/t3/t1/p_1_in [0]),
        .I5(\r7/t3/t1/p_0_in [0]),
        .O(\r7/p_0_out [56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[56]_i_1__6 
       (.I0(\r8/t0/t2/p_0_in [0]),
        .I1(\r8/t2/t0/p_1_in [0]),
        .I2(\r8/t1/t3/p_0_in [0]),
        .I3(k7b[56]),
        .I4(\r8/t3/t1/p_1_in [0]),
        .I5(\r8/t3/t1/p_0_in [0]),
        .O(\r8/p_0_out [56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[56]_i_1__7 
       (.I0(\r9/t0/t2/p_0_in [0]),
        .I1(\r9/t2/t0/p_1_in [0]),
        .I2(\r9/t1/t3/p_0_in [0]),
        .I3(k8b[56]),
        .I4(\r9/t3/t1/p_1_in [0]),
        .I5(\r9/t3/t1/p_0_in [0]),
        .O(\r9/p_0_out [56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair350" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[56]_i_1__8 
       (.I0(\a10/k2a [24]),
        .I1(\a10/k4a [24]),
        .I2(\rf/p_1_in [24]),
        .O(\rf/p_4_out [56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[57]_i_1 
       (.I0(\r1/t0/t2/p_0_in [1]),
        .I1(\r1/t2/t0/p_1_in [1]),
        .I2(\r1/t1/t3/p_0_in [1]),
        .I3(k0b[57]),
        .I4(\r1/t3/t1/p_1_in [1]),
        .I5(\r1/t3/t1/p_0_in [1]),
        .O(\r1/p_0_out [57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[57]_i_1__0 
       (.I0(\r2/t0/t2/p_0_in [1]),
        .I1(\r2/t2/t0/p_1_in [1]),
        .I2(\r2/t1/t3/p_0_in [1]),
        .I3(k1b[57]),
        .I4(\r2/t3/t1/p_1_in [1]),
        .I5(\r2/t3/t1/p_0_in [1]),
        .O(\r2/p_0_out [57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[57]_i_1__1 
       (.I0(\r3/t0/t2/p_0_in [1]),
        .I1(\r3/t2/t0/p_1_in [1]),
        .I2(\r3/t1/t3/p_0_in [1]),
        .I3(k2b[57]),
        .I4(\r3/t3/t1/p_1_in [1]),
        .I5(\r3/t3/t1/p_0_in [1]),
        .O(\r3/p_0_out [57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[57]_i_1__2 
       (.I0(\r4/t0/t2/p_0_in [1]),
        .I1(\r4/t2/t0/p_1_in [1]),
        .I2(\r4/t1/t3/p_0_in [1]),
        .I3(k3b[57]),
        .I4(\r4/t3/t1/p_1_in [1]),
        .I5(\r4/t3/t1/p_0_in [1]),
        .O(\r4/p_0_out [57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[57]_i_1__3 
       (.I0(\r5/t0/t2/p_0_in [1]),
        .I1(\r5/t2/t0/p_1_in [1]),
        .I2(\r5/t1/t3/p_0_in [1]),
        .I3(k4b[57]),
        .I4(\r5/t3/t1/p_1_in [1]),
        .I5(\r5/t3/t1/p_0_in [1]),
        .O(\r5/p_0_out [57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[57]_i_1__4 
       (.I0(\r6/t0/t2/p_0_in [1]),
        .I1(\r6/t2/t0/p_1_in [1]),
        .I2(\r6/t1/t3/p_0_in [1]),
        .I3(k5b[57]),
        .I4(\r6/t3/t1/p_1_in [1]),
        .I5(\r6/t3/t1/p_0_in [1]),
        .O(\r6/p_0_out [57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[57]_i_1__5 
       (.I0(\r7/t0/t2/p_0_in [1]),
        .I1(\r7/t2/t0/p_1_in [1]),
        .I2(\r7/t1/t3/p_0_in [1]),
        .I3(k6b[57]),
        .I4(\r7/t3/t1/p_1_in [1]),
        .I5(\r7/t3/t1/p_0_in [1]),
        .O(\r7/p_0_out [57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[57]_i_1__6 
       (.I0(\r8/t0/t2/p_0_in [1]),
        .I1(\r8/t2/t0/p_1_in [1]),
        .I2(\r8/t1/t3/p_0_in [1]),
        .I3(k7b[57]),
        .I4(\r8/t3/t1/p_1_in [1]),
        .I5(\r8/t3/t1/p_0_in [1]),
        .O(\r8/p_0_out [57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[57]_i_1__7 
       (.I0(\r9/t0/t2/p_0_in [1]),
        .I1(\r9/t2/t0/p_1_in [1]),
        .I2(\r9/t1/t3/p_0_in [1]),
        .I3(k8b[57]),
        .I4(\r9/t3/t1/p_1_in [1]),
        .I5(\r9/t3/t1/p_0_in [1]),
        .O(\r9/p_0_out [57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair349" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[57]_i_1__8 
       (.I0(\a10/k2a [25]),
        .I1(\a10/k4a [25]),
        .I2(\rf/p_1_in [25]),
        .O(\rf/p_4_out [57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[58]_i_1 
       (.I0(\r1/t0/t2/p_0_in [2]),
        .I1(\r1/t2/t0/p_1_in [2]),
        .I2(\r1/t1/t3/p_0_in [2]),
        .I3(k0b[58]),
        .I4(\r1/t3/t1/p_1_in [2]),
        .I5(\r1/t3/t1/p_0_in [2]),
        .O(\r1/p_0_out [58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[58]_i_1__0 
       (.I0(\r2/t0/t2/p_0_in [2]),
        .I1(\r2/t2/t0/p_1_in [2]),
        .I2(\r2/t1/t3/p_0_in [2]),
        .I3(k1b[58]),
        .I4(\r2/t3/t1/p_1_in [2]),
        .I5(\r2/t3/t1/p_0_in [2]),
        .O(\r2/p_0_out [58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[58]_i_1__1 
       (.I0(\r3/t0/t2/p_0_in [2]),
        .I1(\r3/t2/t0/p_1_in [2]),
        .I2(\r3/t1/t3/p_0_in [2]),
        .I3(k2b[58]),
        .I4(\r3/t3/t1/p_1_in [2]),
        .I5(\r3/t3/t1/p_0_in [2]),
        .O(\r3/p_0_out [58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[58]_i_1__2 
       (.I0(\r4/t0/t2/p_0_in [2]),
        .I1(\r4/t2/t0/p_1_in [2]),
        .I2(\r4/t1/t3/p_0_in [2]),
        .I3(k3b[58]),
        .I4(\r4/t3/t1/p_1_in [2]),
        .I5(\r4/t3/t1/p_0_in [2]),
        .O(\r4/p_0_out [58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[58]_i_1__3 
       (.I0(\r5/t0/t2/p_0_in [2]),
        .I1(\r5/t2/t0/p_1_in [2]),
        .I2(\r5/t1/t3/p_0_in [2]),
        .I3(k4b[58]),
        .I4(\r5/t3/t1/p_1_in [2]),
        .I5(\r5/t3/t1/p_0_in [2]),
        .O(\r5/p_0_out [58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[58]_i_1__4 
       (.I0(\r6/t0/t2/p_0_in [2]),
        .I1(\r6/t2/t0/p_1_in [2]),
        .I2(\r6/t1/t3/p_0_in [2]),
        .I3(k5b[58]),
        .I4(\r6/t3/t1/p_1_in [2]),
        .I5(\r6/t3/t1/p_0_in [2]),
        .O(\r6/p_0_out [58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[58]_i_1__5 
       (.I0(\r7/t0/t2/p_0_in [2]),
        .I1(\r7/t2/t0/p_1_in [2]),
        .I2(\r7/t1/t3/p_0_in [2]),
        .I3(k6b[58]),
        .I4(\r7/t3/t1/p_1_in [2]),
        .I5(\r7/t3/t1/p_0_in [2]),
        .O(\r7/p_0_out [58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[58]_i_1__6 
       (.I0(\r8/t0/t2/p_0_in [2]),
        .I1(\r8/t2/t0/p_1_in [2]),
        .I2(\r8/t1/t3/p_0_in [2]),
        .I3(k7b[58]),
        .I4(\r8/t3/t1/p_1_in [2]),
        .I5(\r8/t3/t1/p_0_in [2]),
        .O(\r8/p_0_out [58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[58]_i_1__7 
       (.I0(\r9/t0/t2/p_0_in [2]),
        .I1(\r9/t2/t0/p_1_in [2]),
        .I2(\r9/t1/t3/p_0_in [2]),
        .I3(k8b[58]),
        .I4(\r9/t3/t1/p_1_in [2]),
        .I5(\r9/t3/t1/p_0_in [2]),
        .O(\r9/p_0_out [58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair348" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[58]_i_1__8 
       (.I0(\a10/k2a [26]),
        .I1(\a10/k4a [26]),
        .I2(\rf/p_1_in [26]),
        .O(\rf/p_4_out [58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[59]_i_1 
       (.I0(\r1/t0/t2/p_0_in [3]),
        .I1(\r1/t2/t0/p_1_in [3]),
        .I2(\r1/t1/t3/p_0_in [3]),
        .I3(k0b[59]),
        .I4(\r1/t3/t1/p_1_in [3]),
        .I5(\r1/t3/t1/p_0_in [3]),
        .O(\r1/p_0_out [59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[59]_i_1__0 
       (.I0(\r2/t0/t2/p_0_in [3]),
        .I1(\r2/t2/t0/p_1_in [3]),
        .I2(\r2/t1/t3/p_0_in [3]),
        .I3(k1b[59]),
        .I4(\r2/t3/t1/p_1_in [3]),
        .I5(\r2/t3/t1/p_0_in [3]),
        .O(\r2/p_0_out [59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[59]_i_1__1 
       (.I0(\r3/t0/t2/p_0_in [3]),
        .I1(\r3/t2/t0/p_1_in [3]),
        .I2(\r3/t1/t3/p_0_in [3]),
        .I3(k2b[59]),
        .I4(\r3/t3/t1/p_1_in [3]),
        .I5(\r3/t3/t1/p_0_in [3]),
        .O(\r3/p_0_out [59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[59]_i_1__2 
       (.I0(\r4/t0/t2/p_0_in [3]),
        .I1(\r4/t2/t0/p_1_in [3]),
        .I2(\r4/t1/t3/p_0_in [3]),
        .I3(k3b[59]),
        .I4(\r4/t3/t1/p_1_in [3]),
        .I5(\r4/t3/t1/p_0_in [3]),
        .O(\r4/p_0_out [59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[59]_i_1__3 
       (.I0(\r5/t0/t2/p_0_in [3]),
        .I1(\r5/t2/t0/p_1_in [3]),
        .I2(\r5/t1/t3/p_0_in [3]),
        .I3(k4b[59]),
        .I4(\r5/t3/t1/p_1_in [3]),
        .I5(\r5/t3/t1/p_0_in [3]),
        .O(\r5/p_0_out [59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[59]_i_1__4 
       (.I0(\r6/t0/t2/p_0_in [3]),
        .I1(\r6/t2/t0/p_1_in [3]),
        .I2(\r6/t1/t3/p_0_in [3]),
        .I3(k5b[59]),
        .I4(\r6/t3/t1/p_1_in [3]),
        .I5(\r6/t3/t1/p_0_in [3]),
        .O(\r6/p_0_out [59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[59]_i_1__5 
       (.I0(\r7/t0/t2/p_0_in [3]),
        .I1(\r7/t2/t0/p_1_in [3]),
        .I2(\r7/t1/t3/p_0_in [3]),
        .I3(k6b[59]),
        .I4(\r7/t3/t1/p_1_in [3]),
        .I5(\r7/t3/t1/p_0_in [3]),
        .O(\r7/p_0_out [59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[59]_i_1__6 
       (.I0(\r8/t0/t2/p_0_in [3]),
        .I1(\r8/t2/t0/p_1_in [3]),
        .I2(\r8/t1/t3/p_0_in [3]),
        .I3(k7b[59]),
        .I4(\r8/t3/t1/p_1_in [3]),
        .I5(\r8/t3/t1/p_0_in [3]),
        .O(\r8/p_0_out [59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[59]_i_1__7 
       (.I0(\r9/t0/t2/p_0_in [3]),
        .I1(\r9/t2/t0/p_1_in [3]),
        .I2(\r9/t1/t3/p_0_in [3]),
        .I3(k8b[59]),
        .I4(\r9/t3/t1/p_1_in [3]),
        .I5(\r9/t3/t1/p_0_in [3]),
        .O(\r9/p_0_out [59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair347" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[59]_i_1__8 
       (.I0(\a10/k2a [27]),
        .I1(\a10/k4a [27]),
        .I2(\rf/p_1_in [27]),
        .O(\rf/p_4_out [59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[5]_i_1 
       (.I0(\r1/t0/t1/p_0_in [5]),
        .I1(\r1/t2/t3/p_1_in [5]),
        .I2(\r1/t1/t2/p_0_in [5]),
        .I3(k0b[5]),
        .I4(\r1/t3/t0/p_1_in [5]),
        .I5(\r1/t3/t0/p_0_in [5]),
        .O(\r1/p_0_out [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[5]_i_1__0 
       (.I0(\r2/t0/t1/p_0_in [5]),
        .I1(\r2/t2/t3/p_1_in [5]),
        .I2(\r2/t1/t2/p_0_in [5]),
        .I3(k1b[5]),
        .I4(\r2/t3/t0/p_1_in [5]),
        .I5(\r2/t3/t0/p_0_in [5]),
        .O(\r2/p_0_out [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[5]_i_1__1 
       (.I0(\r3/t0/t1/p_0_in [5]),
        .I1(\r3/t2/t3/p_1_in [5]),
        .I2(\r3/t1/t2/p_0_in [5]),
        .I3(k2b[5]),
        .I4(\r3/t3/t0/p_1_in [5]),
        .I5(\r3/t3/t0/p_0_in [5]),
        .O(\r3/p_0_out [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[5]_i_1__2 
       (.I0(\r4/t0/t1/p_0_in [5]),
        .I1(\r4/t2/t3/p_1_in [5]),
        .I2(\r4/t1/t2/p_0_in [5]),
        .I3(k3b[5]),
        .I4(\r4/t3/t0/p_1_in [5]),
        .I5(\r4/t3/t0/p_0_in [5]),
        .O(\r4/p_0_out [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[5]_i_1__3 
       (.I0(\r5/t0/t1/p_0_in [5]),
        .I1(\r5/t2/t3/p_1_in [5]),
        .I2(\r5/t1/t2/p_0_in [5]),
        .I3(k4b[5]),
        .I4(\r5/t3/t0/p_1_in [5]),
        .I5(\r5/t3/t0/p_0_in [5]),
        .O(\r5/p_0_out [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[5]_i_1__4 
       (.I0(\r6/t0/t1/p_0_in [5]),
        .I1(\r6/t2/t3/p_1_in [5]),
        .I2(\r6/t1/t2/p_0_in [5]),
        .I3(k5b[5]),
        .I4(\r6/t3/t0/p_1_in [5]),
        .I5(\r6/t3/t0/p_0_in [5]),
        .O(\r6/p_0_out [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[5]_i_1__5 
       (.I0(\r7/t0/t1/p_0_in [5]),
        .I1(\r7/t2/t3/p_1_in [5]),
        .I2(\r7/t1/t2/p_0_in [5]),
        .I3(k6b[5]),
        .I4(\r7/t3/t0/p_1_in [5]),
        .I5(\r7/t3/t0/p_0_in [5]),
        .O(\r7/p_0_out [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[5]_i_1__6 
       (.I0(\r8/t0/t1/p_0_in [5]),
        .I1(\r8/t2/t3/p_1_in [5]),
        .I2(\r8/t1/t2/p_0_in [5]),
        .I3(k7b[5]),
        .I4(\r8/t3/t0/p_1_in [5]),
        .I5(\r8/t3/t0/p_0_in [5]),
        .O(\r8/p_0_out [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[5]_i_1__7 
       (.I0(\r9/t0/t1/p_0_in [5]),
        .I1(\r9/t2/t3/p_1_in [5]),
        .I2(\r9/t1/t2/p_0_in [5]),
        .I3(k8b[5]),
        .I4(\r9/t3/t0/p_1_in [5]),
        .I5(\r9/t3/t0/p_0_in [5]),
        .O(\r9/p_0_out [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair337" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[5]_i_1__8 
       (.I0(\a10/k3a [5]),
        .I1(\a10/k4a [5]),
        .I2(\rf/p_0_in [5]),
        .O(\rf/p_4_out [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[60]_i_1 
       (.I0(\r1/t0/t2/p_0_in [4]),
        .I1(\r1/t2/t0/p_1_in [4]),
        .I2(\r1/t1/t3/p_0_in [4]),
        .I3(k0b[60]),
        .I4(\r1/t3/t1/p_1_in [4]),
        .I5(\r1/t3/t1/p_0_in [4]),
        .O(\r1/p_0_out [60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[60]_i_1__0 
       (.I0(\r2/t0/t2/p_0_in [4]),
        .I1(\r2/t2/t0/p_1_in [4]),
        .I2(\r2/t1/t3/p_0_in [4]),
        .I3(k1b[60]),
        .I4(\r2/t3/t1/p_1_in [4]),
        .I5(\r2/t3/t1/p_0_in [4]),
        .O(\r2/p_0_out [60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[60]_i_1__1 
       (.I0(\r3/t0/t2/p_0_in [4]),
        .I1(\r3/t2/t0/p_1_in [4]),
        .I2(\r3/t1/t3/p_0_in [4]),
        .I3(k2b[60]),
        .I4(\r3/t3/t1/p_1_in [4]),
        .I5(\r3/t3/t1/p_0_in [4]),
        .O(\r3/p_0_out [60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[60]_i_1__2 
       (.I0(\r4/t0/t2/p_0_in [4]),
        .I1(\r4/t2/t0/p_1_in [4]),
        .I2(\r4/t1/t3/p_0_in [4]),
        .I3(k3b[60]),
        .I4(\r4/t3/t1/p_1_in [4]),
        .I5(\r4/t3/t1/p_0_in [4]),
        .O(\r4/p_0_out [60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[60]_i_1__3 
       (.I0(\r5/t0/t2/p_0_in [4]),
        .I1(\r5/t2/t0/p_1_in [4]),
        .I2(\r5/t1/t3/p_0_in [4]),
        .I3(k4b[60]),
        .I4(\r5/t3/t1/p_1_in [4]),
        .I5(\r5/t3/t1/p_0_in [4]),
        .O(\r5/p_0_out [60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[60]_i_1__4 
       (.I0(\r6/t0/t2/p_0_in [4]),
        .I1(\r6/t2/t0/p_1_in [4]),
        .I2(\r6/t1/t3/p_0_in [4]),
        .I3(k5b[60]),
        .I4(\r6/t3/t1/p_1_in [4]),
        .I5(\r6/t3/t1/p_0_in [4]),
        .O(\r6/p_0_out [60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[60]_i_1__5 
       (.I0(\r7/t0/t2/p_0_in [4]),
        .I1(\r7/t2/t0/p_1_in [4]),
        .I2(\r7/t1/t3/p_0_in [4]),
        .I3(k6b[60]),
        .I4(\r7/t3/t1/p_1_in [4]),
        .I5(\r7/t3/t1/p_0_in [4]),
        .O(\r7/p_0_out [60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[60]_i_1__6 
       (.I0(\r8/t0/t2/p_0_in [4]),
        .I1(\r8/t2/t0/p_1_in [4]),
        .I2(\r8/t1/t3/p_0_in [4]),
        .I3(k7b[60]),
        .I4(\r8/t3/t1/p_1_in [4]),
        .I5(\r8/t3/t1/p_0_in [4]),
        .O(\r8/p_0_out [60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[60]_i_1__7 
       (.I0(\r9/t0/t2/p_0_in [4]),
        .I1(\r9/t2/t0/p_1_in [4]),
        .I2(\r9/t1/t3/p_0_in [4]),
        .I3(k8b[60]),
        .I4(\r9/t3/t1/p_1_in [4]),
        .I5(\r9/t3/t1/p_0_in [4]),
        .O(\r9/p_0_out [60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair346" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[60]_i_1__8 
       (.I0(\a10/k2a [28]),
        .I1(\a10/k4a [28]),
        .I2(\rf/p_1_in [28]),
        .O(\rf/p_4_out [60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[61]_i_1 
       (.I0(\r1/t0/t2/p_0_in [5]),
        .I1(\r1/t2/t0/p_1_in [5]),
        .I2(\r1/t1/t3/p_0_in [5]),
        .I3(k0b[61]),
        .I4(\r1/t3/t1/p_1_in [5]),
        .I5(\r1/t3/t1/p_0_in [5]),
        .O(\r1/p_0_out [61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[61]_i_1__0 
       (.I0(\r2/t0/t2/p_0_in [5]),
        .I1(\r2/t2/t0/p_1_in [5]),
        .I2(\r2/t1/t3/p_0_in [5]),
        .I3(k1b[61]),
        .I4(\r2/t3/t1/p_1_in [5]),
        .I5(\r2/t3/t1/p_0_in [5]),
        .O(\r2/p_0_out [61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[61]_i_1__1 
       (.I0(\r3/t0/t2/p_0_in [5]),
        .I1(\r3/t2/t0/p_1_in [5]),
        .I2(\r3/t1/t3/p_0_in [5]),
        .I3(k2b[61]),
        .I4(\r3/t3/t1/p_1_in [5]),
        .I5(\r3/t3/t1/p_0_in [5]),
        .O(\r3/p_0_out [61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[61]_i_1__2 
       (.I0(\r4/t0/t2/p_0_in [5]),
        .I1(\r4/t2/t0/p_1_in [5]),
        .I2(\r4/t1/t3/p_0_in [5]),
        .I3(k3b[61]),
        .I4(\r4/t3/t1/p_1_in [5]),
        .I5(\r4/t3/t1/p_0_in [5]),
        .O(\r4/p_0_out [61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[61]_i_1__3 
       (.I0(\r5/t0/t2/p_0_in [5]),
        .I1(\r5/t2/t0/p_1_in [5]),
        .I2(\r5/t1/t3/p_0_in [5]),
        .I3(k4b[61]),
        .I4(\r5/t3/t1/p_1_in [5]),
        .I5(\r5/t3/t1/p_0_in [5]),
        .O(\r5/p_0_out [61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[61]_i_1__4 
       (.I0(\r6/t0/t2/p_0_in [5]),
        .I1(\r6/t2/t0/p_1_in [5]),
        .I2(\r6/t1/t3/p_0_in [5]),
        .I3(k5b[61]),
        .I4(\r6/t3/t1/p_1_in [5]),
        .I5(\r6/t3/t1/p_0_in [5]),
        .O(\r6/p_0_out [61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[61]_i_1__5 
       (.I0(\r7/t0/t2/p_0_in [5]),
        .I1(\r7/t2/t0/p_1_in [5]),
        .I2(\r7/t1/t3/p_0_in [5]),
        .I3(k6b[61]),
        .I4(\r7/t3/t1/p_1_in [5]),
        .I5(\r7/t3/t1/p_0_in [5]),
        .O(\r7/p_0_out [61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[61]_i_1__6 
       (.I0(\r8/t0/t2/p_0_in [5]),
        .I1(\r8/t2/t0/p_1_in [5]),
        .I2(\r8/t1/t3/p_0_in [5]),
        .I3(k7b[61]),
        .I4(\r8/t3/t1/p_1_in [5]),
        .I5(\r8/t3/t1/p_0_in [5]),
        .O(\r8/p_0_out [61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[61]_i_1__7 
       (.I0(\r9/t0/t2/p_0_in [5]),
        .I1(\r9/t2/t0/p_1_in [5]),
        .I2(\r9/t1/t3/p_0_in [5]),
        .I3(k8b[61]),
        .I4(\r9/t3/t1/p_1_in [5]),
        .I5(\r9/t3/t1/p_0_in [5]),
        .O(\r9/p_0_out [61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair345" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[61]_i_1__8 
       (.I0(\a10/k2a [29]),
        .I1(\a10/k4a [29]),
        .I2(\rf/p_1_in [29]),
        .O(\rf/p_4_out [61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[62]_i_1 
       (.I0(\r1/t0/t2/p_0_in [6]),
        .I1(\r1/t2/t0/p_1_in [6]),
        .I2(\r1/t1/t3/p_0_in [6]),
        .I3(k0b[62]),
        .I4(\r1/t3/t1/p_1_in [6]),
        .I5(\r1/t3/t1/p_0_in [6]),
        .O(\r1/p_0_out [62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[62]_i_1__0 
       (.I0(\r2/t0/t2/p_0_in [6]),
        .I1(\r2/t2/t0/p_1_in [6]),
        .I2(\r2/t1/t3/p_0_in [6]),
        .I3(k1b[62]),
        .I4(\r2/t3/t1/p_1_in [6]),
        .I5(\r2/t3/t1/p_0_in [6]),
        .O(\r2/p_0_out [62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[62]_i_1__1 
       (.I0(\r3/t0/t2/p_0_in [6]),
        .I1(\r3/t2/t0/p_1_in [6]),
        .I2(\r3/t1/t3/p_0_in [6]),
        .I3(k2b[62]),
        .I4(\r3/t3/t1/p_1_in [6]),
        .I5(\r3/t3/t1/p_0_in [6]),
        .O(\r3/p_0_out [62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[62]_i_1__2 
       (.I0(\r4/t0/t2/p_0_in [6]),
        .I1(\r4/t2/t0/p_1_in [6]),
        .I2(\r4/t1/t3/p_0_in [6]),
        .I3(k3b[62]),
        .I4(\r4/t3/t1/p_1_in [6]),
        .I5(\r4/t3/t1/p_0_in [6]),
        .O(\r4/p_0_out [62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[62]_i_1__3 
       (.I0(\r5/t0/t2/p_0_in [6]),
        .I1(\r5/t2/t0/p_1_in [6]),
        .I2(\r5/t1/t3/p_0_in [6]),
        .I3(k4b[62]),
        .I4(\r5/t3/t1/p_1_in [6]),
        .I5(\r5/t3/t1/p_0_in [6]),
        .O(\r5/p_0_out [62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[62]_i_1__4 
       (.I0(\r6/t0/t2/p_0_in [6]),
        .I1(\r6/t2/t0/p_1_in [6]),
        .I2(\r6/t1/t3/p_0_in [6]),
        .I3(k5b[62]),
        .I4(\r6/t3/t1/p_1_in [6]),
        .I5(\r6/t3/t1/p_0_in [6]),
        .O(\r6/p_0_out [62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[62]_i_1__5 
       (.I0(\r7/t0/t2/p_0_in [6]),
        .I1(\r7/t2/t0/p_1_in [6]),
        .I2(\r7/t1/t3/p_0_in [6]),
        .I3(k6b[62]),
        .I4(\r7/t3/t1/p_1_in [6]),
        .I5(\r7/t3/t1/p_0_in [6]),
        .O(\r7/p_0_out [62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[62]_i_1__6 
       (.I0(\r8/t0/t2/p_0_in [6]),
        .I1(\r8/t2/t0/p_1_in [6]),
        .I2(\r8/t1/t3/p_0_in [6]),
        .I3(k7b[62]),
        .I4(\r8/t3/t1/p_1_in [6]),
        .I5(\r8/t3/t1/p_0_in [6]),
        .O(\r8/p_0_out [62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[62]_i_1__7 
       (.I0(\r9/t0/t2/p_0_in [6]),
        .I1(\r9/t2/t0/p_1_in [6]),
        .I2(\r9/t1/t3/p_0_in [6]),
        .I3(k8b[62]),
        .I4(\r9/t3/t1/p_1_in [6]),
        .I5(\r9/t3/t1/p_0_in [6]),
        .O(\r9/p_0_out [62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair344" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[62]_i_1__8 
       (.I0(\a10/k2a [30]),
        .I1(\a10/k4a [30]),
        .I2(\rf/p_1_in [30]),
        .O(\rf/p_4_out [62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[63]_i_1 
       (.I0(\r1/t0/t2/p_0_in [7]),
        .I1(\r1/t2/t0/p_1_in [7]),
        .I2(\r1/t1/t3/p_0_in [7]),
        .I3(k0b[63]),
        .I4(\r1/t3/t1/p_1_in [7]),
        .I5(\r1/t3/t1/p_0_in [7]),
        .O(\r1/p_0_out [63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[63]_i_1__0 
       (.I0(\r2/t0/t2/p_0_in [7]),
        .I1(\r2/t2/t0/p_1_in [7]),
        .I2(\r2/t1/t3/p_0_in [7]),
        .I3(k1b[63]),
        .I4(\r2/t3/t1/p_1_in [7]),
        .I5(\r2/t3/t1/p_0_in [7]),
        .O(\r2/p_0_out [63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[63]_i_1__1 
       (.I0(\r3/t0/t2/p_0_in [7]),
        .I1(\r3/t2/t0/p_1_in [7]),
        .I2(\r3/t1/t3/p_0_in [7]),
        .I3(k2b[63]),
        .I4(\r3/t3/t1/p_1_in [7]),
        .I5(\r3/t3/t1/p_0_in [7]),
        .O(\r3/p_0_out [63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[63]_i_1__2 
       (.I0(\r4/t0/t2/p_0_in [7]),
        .I1(\r4/t2/t0/p_1_in [7]),
        .I2(\r4/t1/t3/p_0_in [7]),
        .I3(k3b[63]),
        .I4(\r4/t3/t1/p_1_in [7]),
        .I5(\r4/t3/t1/p_0_in [7]),
        .O(\r4/p_0_out [63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[63]_i_1__3 
       (.I0(\r5/t0/t2/p_0_in [7]),
        .I1(\r5/t2/t0/p_1_in [7]),
        .I2(\r5/t1/t3/p_0_in [7]),
        .I3(k4b[63]),
        .I4(\r5/t3/t1/p_1_in [7]),
        .I5(\r5/t3/t1/p_0_in [7]),
        .O(\r5/p_0_out [63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[63]_i_1__4 
       (.I0(\r6/t0/t2/p_0_in [7]),
        .I1(\r6/t2/t0/p_1_in [7]),
        .I2(\r6/t1/t3/p_0_in [7]),
        .I3(k5b[63]),
        .I4(\r6/t3/t1/p_1_in [7]),
        .I5(\r6/t3/t1/p_0_in [7]),
        .O(\r6/p_0_out [63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[63]_i_1__5 
       (.I0(\r7/t0/t2/p_0_in [7]),
        .I1(\r7/t2/t0/p_1_in [7]),
        .I2(\r7/t1/t3/p_0_in [7]),
        .I3(k6b[63]),
        .I4(\r7/t3/t1/p_1_in [7]),
        .I5(\r7/t3/t1/p_0_in [7]),
        .O(\r7/p_0_out [63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[63]_i_1__6 
       (.I0(\r8/t0/t2/p_0_in [7]),
        .I1(\r8/t2/t0/p_1_in [7]),
        .I2(\r8/t1/t3/p_0_in [7]),
        .I3(k7b[63]),
        .I4(\r8/t3/t1/p_1_in [7]),
        .I5(\r8/t3/t1/p_0_in [7]),
        .O(\r8/p_0_out [63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[63]_i_1__7 
       (.I0(\r9/t0/t2/p_0_in [7]),
        .I1(\r9/t2/t0/p_1_in [7]),
        .I2(\r9/t1/t3/p_0_in [7]),
        .I3(k8b[63]),
        .I4(\r9/t3/t1/p_1_in [7]),
        .I5(\r9/t3/t1/p_0_in [7]),
        .O(\r9/p_0_out [63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair343" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[63]_i_1__8 
       (.I0(\a10/k2a [31]),
        .I1(\a10/k4a [31]),
        .I2(\rf/p_1_in [31]),
        .O(\rf/p_4_out [63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[64]_i_1 
       (.I0(\r1/t0/t3/p_1_in [0]),
        .I1(\r1/t2/t1/p_0_in [0]),
        .I2(\r1/t1/t0/p_1_in [0]),
        .I3(\r1/t1/t0/p_0_in [0]),
        .I4(k0b[64]),
        .I5(\r1/t3/t2/p_0_in [0]),
        .O(\r1/p_0_out [64]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[64]_i_1__0 
       (.I0(\r2/t0/t3/p_1_in [0]),
        .I1(\r2/t2/t1/p_0_in [0]),
        .I2(\r2/t1/t0/p_1_in [0]),
        .I3(\r2/t1/t0/p_0_in [0]),
        .I4(k1b[64]),
        .I5(\r2/t3/t2/p_0_in [0]),
        .O(\r2/p_0_out [64]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[64]_i_1__1 
       (.I0(\r3/t0/t3/p_1_in [0]),
        .I1(\r3/t2/t1/p_0_in [0]),
        .I2(\r3/t1/t0/p_1_in [0]),
        .I3(\r3/t1/t0/p_0_in [0]),
        .I4(k2b[64]),
        .I5(\r3/t3/t2/p_0_in [0]),
        .O(\r3/p_0_out [64]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[64]_i_1__2 
       (.I0(\r4/t0/t3/p_1_in [0]),
        .I1(\r4/t2/t1/p_0_in [0]),
        .I2(\r4/t1/t0/p_1_in [0]),
        .I3(\r4/t1/t0/p_0_in [0]),
        .I4(k3b[64]),
        .I5(\r4/t3/t2/p_0_in [0]),
        .O(\r4/p_0_out [64]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[64]_i_1__3 
       (.I0(\r5/t0/t3/p_1_in [0]),
        .I1(\r5/t2/t1/p_0_in [0]),
        .I2(\r5/t1/t0/p_1_in [0]),
        .I3(\r5/t1/t0/p_0_in [0]),
        .I4(k4b[64]),
        .I5(\r5/t3/t2/p_0_in [0]),
        .O(\r5/p_0_out [64]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[64]_i_1__4 
       (.I0(\r6/t0/t3/p_1_in [0]),
        .I1(\r6/t2/t1/p_0_in [0]),
        .I2(\r6/t1/t0/p_1_in [0]),
        .I3(\r6/t1/t0/p_0_in [0]),
        .I4(k5b[64]),
        .I5(\r6/t3/t2/p_0_in [0]),
        .O(\r6/p_0_out [64]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[64]_i_1__5 
       (.I0(\r7/t0/t3/p_1_in [0]),
        .I1(\r7/t2/t1/p_0_in [0]),
        .I2(\r7/t1/t0/p_1_in [0]),
        .I3(\r7/t1/t0/p_0_in [0]),
        .I4(k6b[64]),
        .I5(\r7/t3/t2/p_0_in [0]),
        .O(\r7/p_0_out [64]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[64]_i_1__6 
       (.I0(\r8/t0/t3/p_1_in [0]),
        .I1(\r8/t2/t1/p_0_in [0]),
        .I2(\r8/t1/t0/p_1_in [0]),
        .I3(\r8/t1/t0/p_0_in [0]),
        .I4(k7b[64]),
        .I5(\r8/t3/t2/p_0_in [0]),
        .O(\r8/p_0_out [64]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[64]_i_1__7 
       (.I0(\r9/t0/t3/p_1_in [0]),
        .I1(\r9/t2/t1/p_0_in [0]),
        .I2(\r9/t1/t0/p_1_in [0]),
        .I3(\r9/t1/t0/p_0_in [0]),
        .I4(k8b[64]),
        .I5(\r9/t3/t2/p_0_in [0]),
        .O(\r9/p_0_out [64]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair374" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[64]_i_1__8 
       (.I0(\a10/k1a [0]),
        .I1(\a10/k4a [0]),
        .I2(\rf/p_2_in [0]),
        .O(\rf/p_4_out [64]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[65]_i_1 
       (.I0(\r1/t0/t3/p_1_in [1]),
        .I1(\r1/t2/t1/p_0_in [1]),
        .I2(\r1/t1/t0/p_1_in [1]),
        .I3(\r1/t1/t0/p_0_in [1]),
        .I4(k0b[65]),
        .I5(\r1/t3/t2/p_0_in [1]),
        .O(\r1/p_0_out [65]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[65]_i_1__0 
       (.I0(\r2/t0/t3/p_1_in [1]),
        .I1(\r2/t2/t1/p_0_in [1]),
        .I2(\r2/t1/t0/p_1_in [1]),
        .I3(\r2/t1/t0/p_0_in [1]),
        .I4(k1b[65]),
        .I5(\r2/t3/t2/p_0_in [1]),
        .O(\r2/p_0_out [65]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[65]_i_1__1 
       (.I0(\r3/t0/t3/p_1_in [1]),
        .I1(\r3/t2/t1/p_0_in [1]),
        .I2(\r3/t1/t0/p_1_in [1]),
        .I3(\r3/t1/t0/p_0_in [1]),
        .I4(k2b[65]),
        .I5(\r3/t3/t2/p_0_in [1]),
        .O(\r3/p_0_out [65]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[65]_i_1__2 
       (.I0(\r4/t0/t3/p_1_in [1]),
        .I1(\r4/t2/t1/p_0_in [1]),
        .I2(\r4/t1/t0/p_1_in [1]),
        .I3(\r4/t1/t0/p_0_in [1]),
        .I4(k3b[65]),
        .I5(\r4/t3/t2/p_0_in [1]),
        .O(\r4/p_0_out [65]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[65]_i_1__3 
       (.I0(\r5/t0/t3/p_1_in [1]),
        .I1(\r5/t2/t1/p_0_in [1]),
        .I2(\r5/t1/t0/p_1_in [1]),
        .I3(\r5/t1/t0/p_0_in [1]),
        .I4(k4b[65]),
        .I5(\r5/t3/t2/p_0_in [1]),
        .O(\r5/p_0_out [65]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[65]_i_1__4 
       (.I0(\r6/t0/t3/p_1_in [1]),
        .I1(\r6/t2/t1/p_0_in [1]),
        .I2(\r6/t1/t0/p_1_in [1]),
        .I3(\r6/t1/t0/p_0_in [1]),
        .I4(k5b[65]),
        .I5(\r6/t3/t2/p_0_in [1]),
        .O(\r6/p_0_out [65]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[65]_i_1__5 
       (.I0(\r7/t0/t3/p_1_in [1]),
        .I1(\r7/t2/t1/p_0_in [1]),
        .I2(\r7/t1/t0/p_1_in [1]),
        .I3(\r7/t1/t0/p_0_in [1]),
        .I4(k6b[65]),
        .I5(\r7/t3/t2/p_0_in [1]),
        .O(\r7/p_0_out [65]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[65]_i_1__6 
       (.I0(\r8/t0/t3/p_1_in [1]),
        .I1(\r8/t2/t1/p_0_in [1]),
        .I2(\r8/t1/t0/p_1_in [1]),
        .I3(\r8/t1/t0/p_0_in [1]),
        .I4(k7b[65]),
        .I5(\r8/t3/t2/p_0_in [1]),
        .O(\r8/p_0_out [65]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[65]_i_1__7 
       (.I0(\r9/t0/t3/p_1_in [1]),
        .I1(\r9/t2/t1/p_0_in [1]),
        .I2(\r9/t1/t0/p_1_in [1]),
        .I3(\r9/t1/t0/p_0_in [1]),
        .I4(k8b[65]),
        .I5(\r9/t3/t2/p_0_in [1]),
        .O(\r9/p_0_out [65]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair373" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[65]_i_1__8 
       (.I0(\a10/k1a [1]),
        .I1(\a10/k4a [1]),
        .I2(\rf/p_2_in [1]),
        .O(\rf/p_4_out [65]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[66]_i_1 
       (.I0(\r1/t0/t3/p_1_in [2]),
        .I1(\r1/t2/t1/p_0_in [2]),
        .I2(\r1/t1/t0/p_1_in [2]),
        .I3(\r1/t1/t0/p_0_in [2]),
        .I4(k0b[66]),
        .I5(\r1/t3/t2/p_0_in [2]),
        .O(\r1/p_0_out [66]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[66]_i_1__0 
       (.I0(\r2/t0/t3/p_1_in [2]),
        .I1(\r2/t2/t1/p_0_in [2]),
        .I2(\r2/t1/t0/p_1_in [2]),
        .I3(\r2/t1/t0/p_0_in [2]),
        .I4(k1b[66]),
        .I5(\r2/t3/t2/p_0_in [2]),
        .O(\r2/p_0_out [66]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[66]_i_1__1 
       (.I0(\r3/t0/t3/p_1_in [2]),
        .I1(\r3/t2/t1/p_0_in [2]),
        .I2(\r3/t1/t0/p_1_in [2]),
        .I3(\r3/t1/t0/p_0_in [2]),
        .I4(k2b[66]),
        .I5(\r3/t3/t2/p_0_in [2]),
        .O(\r3/p_0_out [66]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[66]_i_1__2 
       (.I0(\r4/t0/t3/p_1_in [2]),
        .I1(\r4/t2/t1/p_0_in [2]),
        .I2(\r4/t1/t0/p_1_in [2]),
        .I3(\r4/t1/t0/p_0_in [2]),
        .I4(k3b[66]),
        .I5(\r4/t3/t2/p_0_in [2]),
        .O(\r4/p_0_out [66]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[66]_i_1__3 
       (.I0(\r5/t0/t3/p_1_in [2]),
        .I1(\r5/t2/t1/p_0_in [2]),
        .I2(\r5/t1/t0/p_1_in [2]),
        .I3(\r5/t1/t0/p_0_in [2]),
        .I4(k4b[66]),
        .I5(\r5/t3/t2/p_0_in [2]),
        .O(\r5/p_0_out [66]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[66]_i_1__4 
       (.I0(\r6/t0/t3/p_1_in [2]),
        .I1(\r6/t2/t1/p_0_in [2]),
        .I2(\r6/t1/t0/p_1_in [2]),
        .I3(\r6/t1/t0/p_0_in [2]),
        .I4(k5b[66]),
        .I5(\r6/t3/t2/p_0_in [2]),
        .O(\r6/p_0_out [66]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[66]_i_1__5 
       (.I0(\r7/t0/t3/p_1_in [2]),
        .I1(\r7/t2/t1/p_0_in [2]),
        .I2(\r7/t1/t0/p_1_in [2]),
        .I3(\r7/t1/t0/p_0_in [2]),
        .I4(k6b[66]),
        .I5(\r7/t3/t2/p_0_in [2]),
        .O(\r7/p_0_out [66]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[66]_i_1__6 
       (.I0(\r8/t0/t3/p_1_in [2]),
        .I1(\r8/t2/t1/p_0_in [2]),
        .I2(\r8/t1/t0/p_1_in [2]),
        .I3(\r8/t1/t0/p_0_in [2]),
        .I4(k7b[66]),
        .I5(\r8/t3/t2/p_0_in [2]),
        .O(\r8/p_0_out [66]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[66]_i_1__7 
       (.I0(\r9/t0/t3/p_1_in [2]),
        .I1(\r9/t2/t1/p_0_in [2]),
        .I2(\r9/t1/t0/p_1_in [2]),
        .I3(\r9/t1/t0/p_0_in [2]),
        .I4(k8b[66]),
        .I5(\r9/t3/t2/p_0_in [2]),
        .O(\r9/p_0_out [66]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair372" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[66]_i_1__8 
       (.I0(\a10/k1a [2]),
        .I1(\a10/k4a [2]),
        .I2(\rf/p_2_in [2]),
        .O(\rf/p_4_out [66]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[67]_i_1 
       (.I0(\r1/t0/t3/p_1_in [3]),
        .I1(\r1/t2/t1/p_0_in [3]),
        .I2(\r1/t1/t0/p_1_in [3]),
        .I3(\r1/t1/t0/p_0_in [3]),
        .I4(k0b[67]),
        .I5(\r1/t3/t2/p_0_in [3]),
        .O(\r1/p_0_out [67]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[67]_i_1__0 
       (.I0(\r2/t0/t3/p_1_in [3]),
        .I1(\r2/t2/t1/p_0_in [3]),
        .I2(\r2/t1/t0/p_1_in [3]),
        .I3(\r2/t1/t0/p_0_in [3]),
        .I4(k1b[67]),
        .I5(\r2/t3/t2/p_0_in [3]),
        .O(\r2/p_0_out [67]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[67]_i_1__1 
       (.I0(\r3/t0/t3/p_1_in [3]),
        .I1(\r3/t2/t1/p_0_in [3]),
        .I2(\r3/t1/t0/p_1_in [3]),
        .I3(\r3/t1/t0/p_0_in [3]),
        .I4(k2b[67]),
        .I5(\r3/t3/t2/p_0_in [3]),
        .O(\r3/p_0_out [67]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[67]_i_1__2 
       (.I0(\r4/t0/t3/p_1_in [3]),
        .I1(\r4/t2/t1/p_0_in [3]),
        .I2(\r4/t1/t0/p_1_in [3]),
        .I3(\r4/t1/t0/p_0_in [3]),
        .I4(k3b[67]),
        .I5(\r4/t3/t2/p_0_in [3]),
        .O(\r4/p_0_out [67]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[67]_i_1__3 
       (.I0(\r5/t0/t3/p_1_in [3]),
        .I1(\r5/t2/t1/p_0_in [3]),
        .I2(\r5/t1/t0/p_1_in [3]),
        .I3(\r5/t1/t0/p_0_in [3]),
        .I4(k4b[67]),
        .I5(\r5/t3/t2/p_0_in [3]),
        .O(\r5/p_0_out [67]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[67]_i_1__4 
       (.I0(\r6/t0/t3/p_1_in [3]),
        .I1(\r6/t2/t1/p_0_in [3]),
        .I2(\r6/t1/t0/p_1_in [3]),
        .I3(\r6/t1/t0/p_0_in [3]),
        .I4(k5b[67]),
        .I5(\r6/t3/t2/p_0_in [3]),
        .O(\r6/p_0_out [67]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[67]_i_1__5 
       (.I0(\r7/t0/t3/p_1_in [3]),
        .I1(\r7/t2/t1/p_0_in [3]),
        .I2(\r7/t1/t0/p_1_in [3]),
        .I3(\r7/t1/t0/p_0_in [3]),
        .I4(k6b[67]),
        .I5(\r7/t3/t2/p_0_in [3]),
        .O(\r7/p_0_out [67]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[67]_i_1__6 
       (.I0(\r8/t0/t3/p_1_in [3]),
        .I1(\r8/t2/t1/p_0_in [3]),
        .I2(\r8/t1/t0/p_1_in [3]),
        .I3(\r8/t1/t0/p_0_in [3]),
        .I4(k7b[67]),
        .I5(\r8/t3/t2/p_0_in [3]),
        .O(\r8/p_0_out [67]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[67]_i_1__7 
       (.I0(\r9/t0/t3/p_1_in [3]),
        .I1(\r9/t2/t1/p_0_in [3]),
        .I2(\r9/t1/t0/p_1_in [3]),
        .I3(\r9/t1/t0/p_0_in [3]),
        .I4(k8b[67]),
        .I5(\r9/t3/t2/p_0_in [3]),
        .O(\r9/p_0_out [67]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair371" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[67]_i_1__8 
       (.I0(\a10/k1a [3]),
        .I1(\a10/k4a [3]),
        .I2(\rf/p_2_in [3]),
        .O(\rf/p_4_out [67]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[68]_i_1 
       (.I0(\r1/t0/t3/p_1_in [4]),
        .I1(\r1/t2/t1/p_0_in [4]),
        .I2(\r1/t1/t0/p_1_in [4]),
        .I3(\r1/t1/t0/p_0_in [4]),
        .I4(k0b[68]),
        .I5(\r1/t3/t2/p_0_in [4]),
        .O(\r1/p_0_out [68]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[68]_i_1__0 
       (.I0(\r2/t0/t3/p_1_in [4]),
        .I1(\r2/t2/t1/p_0_in [4]),
        .I2(\r2/t1/t0/p_1_in [4]),
        .I3(\r2/t1/t0/p_0_in [4]),
        .I4(k1b[68]),
        .I5(\r2/t3/t2/p_0_in [4]),
        .O(\r2/p_0_out [68]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[68]_i_1__1 
       (.I0(\r3/t0/t3/p_1_in [4]),
        .I1(\r3/t2/t1/p_0_in [4]),
        .I2(\r3/t1/t0/p_1_in [4]),
        .I3(\r3/t1/t0/p_0_in [4]),
        .I4(k2b[68]),
        .I5(\r3/t3/t2/p_0_in [4]),
        .O(\r3/p_0_out [68]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[68]_i_1__2 
       (.I0(\r4/t0/t3/p_1_in [4]),
        .I1(\r4/t2/t1/p_0_in [4]),
        .I2(\r4/t1/t0/p_1_in [4]),
        .I3(\r4/t1/t0/p_0_in [4]),
        .I4(k3b[68]),
        .I5(\r4/t3/t2/p_0_in [4]),
        .O(\r4/p_0_out [68]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[68]_i_1__3 
       (.I0(\r5/t0/t3/p_1_in [4]),
        .I1(\r5/t2/t1/p_0_in [4]),
        .I2(\r5/t1/t0/p_1_in [4]),
        .I3(\r5/t1/t0/p_0_in [4]),
        .I4(k4b[68]),
        .I5(\r5/t3/t2/p_0_in [4]),
        .O(\r5/p_0_out [68]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[68]_i_1__4 
       (.I0(\r6/t0/t3/p_1_in [4]),
        .I1(\r6/t2/t1/p_0_in [4]),
        .I2(\r6/t1/t0/p_1_in [4]),
        .I3(\r6/t1/t0/p_0_in [4]),
        .I4(k5b[68]),
        .I5(\r6/t3/t2/p_0_in [4]),
        .O(\r6/p_0_out [68]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[68]_i_1__5 
       (.I0(\r7/t0/t3/p_1_in [4]),
        .I1(\r7/t2/t1/p_0_in [4]),
        .I2(\r7/t1/t0/p_1_in [4]),
        .I3(\r7/t1/t0/p_0_in [4]),
        .I4(k6b[68]),
        .I5(\r7/t3/t2/p_0_in [4]),
        .O(\r7/p_0_out [68]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[68]_i_1__6 
       (.I0(\r8/t0/t3/p_1_in [4]),
        .I1(\r8/t2/t1/p_0_in [4]),
        .I2(\r8/t1/t0/p_1_in [4]),
        .I3(\r8/t1/t0/p_0_in [4]),
        .I4(k7b[68]),
        .I5(\r8/t3/t2/p_0_in [4]),
        .O(\r8/p_0_out [68]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[68]_i_1__7 
       (.I0(\r9/t0/t3/p_1_in [4]),
        .I1(\r9/t2/t1/p_0_in [4]),
        .I2(\r9/t1/t0/p_1_in [4]),
        .I3(\r9/t1/t0/p_0_in [4]),
        .I4(k8b[68]),
        .I5(\r9/t3/t2/p_0_in [4]),
        .O(\r9/p_0_out [68]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair370" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[68]_i_1__8 
       (.I0(\a10/k1a [4]),
        .I1(\a10/k4a [4]),
        .I2(\rf/p_2_in [4]),
        .O(\rf/p_4_out [68]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[69]_i_1 
       (.I0(\r1/t0/t3/p_1_in [5]),
        .I1(\r1/t2/t1/p_0_in [5]),
        .I2(\r1/t1/t0/p_1_in [5]),
        .I3(\r1/t1/t0/p_0_in [5]),
        .I4(k0b[69]),
        .I5(\r1/t3/t2/p_0_in [5]),
        .O(\r1/p_0_out [69]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[69]_i_1__0 
       (.I0(\r2/t0/t3/p_1_in [5]),
        .I1(\r2/t2/t1/p_0_in [5]),
        .I2(\r2/t1/t0/p_1_in [5]),
        .I3(\r2/t1/t0/p_0_in [5]),
        .I4(k1b[69]),
        .I5(\r2/t3/t2/p_0_in [5]),
        .O(\r2/p_0_out [69]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[69]_i_1__1 
       (.I0(\r3/t0/t3/p_1_in [5]),
        .I1(\r3/t2/t1/p_0_in [5]),
        .I2(\r3/t1/t0/p_1_in [5]),
        .I3(\r3/t1/t0/p_0_in [5]),
        .I4(k2b[69]),
        .I5(\r3/t3/t2/p_0_in [5]),
        .O(\r3/p_0_out [69]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[69]_i_1__2 
       (.I0(\r4/t0/t3/p_1_in [5]),
        .I1(\r4/t2/t1/p_0_in [5]),
        .I2(\r4/t1/t0/p_1_in [5]),
        .I3(\r4/t1/t0/p_0_in [5]),
        .I4(k3b[69]),
        .I5(\r4/t3/t2/p_0_in [5]),
        .O(\r4/p_0_out [69]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[69]_i_1__3 
       (.I0(\r5/t0/t3/p_1_in [5]),
        .I1(\r5/t2/t1/p_0_in [5]),
        .I2(\r5/t1/t0/p_1_in [5]),
        .I3(\r5/t1/t0/p_0_in [5]),
        .I4(k4b[69]),
        .I5(\r5/t3/t2/p_0_in [5]),
        .O(\r5/p_0_out [69]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[69]_i_1__4 
       (.I0(\r6/t0/t3/p_1_in [5]),
        .I1(\r6/t2/t1/p_0_in [5]),
        .I2(\r6/t1/t0/p_1_in [5]),
        .I3(\r6/t1/t0/p_0_in [5]),
        .I4(k5b[69]),
        .I5(\r6/t3/t2/p_0_in [5]),
        .O(\r6/p_0_out [69]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[69]_i_1__5 
       (.I0(\r7/t0/t3/p_1_in [5]),
        .I1(\r7/t2/t1/p_0_in [5]),
        .I2(\r7/t1/t0/p_1_in [5]),
        .I3(\r7/t1/t0/p_0_in [5]),
        .I4(k6b[69]),
        .I5(\r7/t3/t2/p_0_in [5]),
        .O(\r7/p_0_out [69]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[69]_i_1__6 
       (.I0(\r8/t0/t3/p_1_in [5]),
        .I1(\r8/t2/t1/p_0_in [5]),
        .I2(\r8/t1/t0/p_1_in [5]),
        .I3(\r8/t1/t0/p_0_in [5]),
        .I4(k7b[69]),
        .I5(\r8/t3/t2/p_0_in [5]),
        .O(\r8/p_0_out [69]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[69]_i_1__7 
       (.I0(\r9/t0/t3/p_1_in [5]),
        .I1(\r9/t2/t1/p_0_in [5]),
        .I2(\r9/t1/t0/p_1_in [5]),
        .I3(\r9/t1/t0/p_0_in [5]),
        .I4(k8b[69]),
        .I5(\r9/t3/t2/p_0_in [5]),
        .O(\r9/p_0_out [69]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair369" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[69]_i_1__8 
       (.I0(\a10/k1a [5]),
        .I1(\a10/k4a [5]),
        .I2(\rf/p_2_in [5]),
        .O(\rf/p_4_out [69]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[6]_i_1 
       (.I0(\r1/t0/t1/p_0_in [6]),
        .I1(\r1/t2/t3/p_1_in [6]),
        .I2(\r1/t1/t2/p_0_in [6]),
        .I3(k0b[6]),
        .I4(\r1/t3/t0/p_1_in [6]),
        .I5(\r1/t3/t0/p_0_in [6]),
        .O(\r1/p_0_out [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[6]_i_1__0 
       (.I0(\r2/t0/t1/p_0_in [6]),
        .I1(\r2/t2/t3/p_1_in [6]),
        .I2(\r2/t1/t2/p_0_in [6]),
        .I3(k1b[6]),
        .I4(\r2/t3/t0/p_1_in [6]),
        .I5(\r2/t3/t0/p_0_in [6]),
        .O(\r2/p_0_out [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[6]_i_1__1 
       (.I0(\r3/t0/t1/p_0_in [6]),
        .I1(\r3/t2/t3/p_1_in [6]),
        .I2(\r3/t1/t2/p_0_in [6]),
        .I3(k2b[6]),
        .I4(\r3/t3/t0/p_1_in [6]),
        .I5(\r3/t3/t0/p_0_in [6]),
        .O(\r3/p_0_out [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[6]_i_1__2 
       (.I0(\r4/t0/t1/p_0_in [6]),
        .I1(\r4/t2/t3/p_1_in [6]),
        .I2(\r4/t1/t2/p_0_in [6]),
        .I3(k3b[6]),
        .I4(\r4/t3/t0/p_1_in [6]),
        .I5(\r4/t3/t0/p_0_in [6]),
        .O(\r4/p_0_out [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[6]_i_1__3 
       (.I0(\r5/t0/t1/p_0_in [6]),
        .I1(\r5/t2/t3/p_1_in [6]),
        .I2(\r5/t1/t2/p_0_in [6]),
        .I3(k4b[6]),
        .I4(\r5/t3/t0/p_1_in [6]),
        .I5(\r5/t3/t0/p_0_in [6]),
        .O(\r5/p_0_out [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[6]_i_1__4 
       (.I0(\r6/t0/t1/p_0_in [6]),
        .I1(\r6/t2/t3/p_1_in [6]),
        .I2(\r6/t1/t2/p_0_in [6]),
        .I3(k5b[6]),
        .I4(\r6/t3/t0/p_1_in [6]),
        .I5(\r6/t3/t0/p_0_in [6]),
        .O(\r6/p_0_out [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[6]_i_1__5 
       (.I0(\r7/t0/t1/p_0_in [6]),
        .I1(\r7/t2/t3/p_1_in [6]),
        .I2(\r7/t1/t2/p_0_in [6]),
        .I3(k6b[6]),
        .I4(\r7/t3/t0/p_1_in [6]),
        .I5(\r7/t3/t0/p_0_in [6]),
        .O(\r7/p_0_out [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[6]_i_1__6 
       (.I0(\r8/t0/t1/p_0_in [6]),
        .I1(\r8/t2/t3/p_1_in [6]),
        .I2(\r8/t1/t2/p_0_in [6]),
        .I3(k7b[6]),
        .I4(\r8/t3/t0/p_1_in [6]),
        .I5(\r8/t3/t0/p_0_in [6]),
        .O(\r8/p_0_out [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[6]_i_1__7 
       (.I0(\r9/t0/t1/p_0_in [6]),
        .I1(\r9/t2/t3/p_1_in [6]),
        .I2(\r9/t1/t2/p_0_in [6]),
        .I3(k8b[6]),
        .I4(\r9/t3/t0/p_1_in [6]),
        .I5(\r9/t3/t0/p_0_in [6]),
        .O(\r9/p_0_out [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair336" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[6]_i_1__8 
       (.I0(\a10/k3a [6]),
        .I1(\a10/k4a [6]),
        .I2(\rf/p_0_in [6]),
        .O(\rf/p_4_out [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[70]_i_1 
       (.I0(\r1/t0/t3/p_1_in [6]),
        .I1(\r1/t2/t1/p_0_in [6]),
        .I2(\r1/t1/t0/p_1_in [6]),
        .I3(\r1/t1/t0/p_0_in [6]),
        .I4(k0b[70]),
        .I5(\r1/t3/t2/p_0_in [6]),
        .O(\r1/p_0_out [70]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[70]_i_1__0 
       (.I0(\r2/t0/t3/p_1_in [6]),
        .I1(\r2/t2/t1/p_0_in [6]),
        .I2(\r2/t1/t0/p_1_in [6]),
        .I3(\r2/t1/t0/p_0_in [6]),
        .I4(k1b[70]),
        .I5(\r2/t3/t2/p_0_in [6]),
        .O(\r2/p_0_out [70]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[70]_i_1__1 
       (.I0(\r3/t0/t3/p_1_in [6]),
        .I1(\r3/t2/t1/p_0_in [6]),
        .I2(\r3/t1/t0/p_1_in [6]),
        .I3(\r3/t1/t0/p_0_in [6]),
        .I4(k2b[70]),
        .I5(\r3/t3/t2/p_0_in [6]),
        .O(\r3/p_0_out [70]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[70]_i_1__2 
       (.I0(\r4/t0/t3/p_1_in [6]),
        .I1(\r4/t2/t1/p_0_in [6]),
        .I2(\r4/t1/t0/p_1_in [6]),
        .I3(\r4/t1/t0/p_0_in [6]),
        .I4(k3b[70]),
        .I5(\r4/t3/t2/p_0_in [6]),
        .O(\r4/p_0_out [70]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[70]_i_1__3 
       (.I0(\r5/t0/t3/p_1_in [6]),
        .I1(\r5/t2/t1/p_0_in [6]),
        .I2(\r5/t1/t0/p_1_in [6]),
        .I3(\r5/t1/t0/p_0_in [6]),
        .I4(k4b[70]),
        .I5(\r5/t3/t2/p_0_in [6]),
        .O(\r5/p_0_out [70]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[70]_i_1__4 
       (.I0(\r6/t0/t3/p_1_in [6]),
        .I1(\r6/t2/t1/p_0_in [6]),
        .I2(\r6/t1/t0/p_1_in [6]),
        .I3(\r6/t1/t0/p_0_in [6]),
        .I4(k5b[70]),
        .I5(\r6/t3/t2/p_0_in [6]),
        .O(\r6/p_0_out [70]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[70]_i_1__5 
       (.I0(\r7/t0/t3/p_1_in [6]),
        .I1(\r7/t2/t1/p_0_in [6]),
        .I2(\r7/t1/t0/p_1_in [6]),
        .I3(\r7/t1/t0/p_0_in [6]),
        .I4(k6b[70]),
        .I5(\r7/t3/t2/p_0_in [6]),
        .O(\r7/p_0_out [70]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[70]_i_1__6 
       (.I0(\r8/t0/t3/p_1_in [6]),
        .I1(\r8/t2/t1/p_0_in [6]),
        .I2(\r8/t1/t0/p_1_in [6]),
        .I3(\r8/t1/t0/p_0_in [6]),
        .I4(k7b[70]),
        .I5(\r8/t3/t2/p_0_in [6]),
        .O(\r8/p_0_out [70]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[70]_i_1__7 
       (.I0(\r9/t0/t3/p_1_in [6]),
        .I1(\r9/t2/t1/p_0_in [6]),
        .I2(\r9/t1/t0/p_1_in [6]),
        .I3(\r9/t1/t0/p_0_in [6]),
        .I4(k8b[70]),
        .I5(\r9/t3/t2/p_0_in [6]),
        .O(\r9/p_0_out [70]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair368" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[70]_i_1__8 
       (.I0(\a10/k1a [6]),
        .I1(\a10/k4a [6]),
        .I2(\rf/p_2_in [6]),
        .O(\rf/p_4_out [70]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[71]_i_1 
       (.I0(\r1/t0/t3/p_1_in [7]),
        .I1(\r1/t2/t1/p_0_in [7]),
        .I2(\r1/t1/t0/p_1_in [7]),
        .I3(\r1/t1/t0/p_0_in [7]),
        .I4(k0b[71]),
        .I5(\r1/t3/t2/p_0_in [7]),
        .O(\r1/p_0_out [71]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[71]_i_1__0 
       (.I0(\r2/t0/t3/p_1_in [7]),
        .I1(\r2/t2/t1/p_0_in [7]),
        .I2(\r2/t1/t0/p_1_in [7]),
        .I3(\r2/t1/t0/p_0_in [7]),
        .I4(k1b[71]),
        .I5(\r2/t3/t2/p_0_in [7]),
        .O(\r2/p_0_out [71]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[71]_i_1__1 
       (.I0(\r3/t0/t3/p_1_in [7]),
        .I1(\r3/t2/t1/p_0_in [7]),
        .I2(\r3/t1/t0/p_1_in [7]),
        .I3(\r3/t1/t0/p_0_in [7]),
        .I4(k2b[71]),
        .I5(\r3/t3/t2/p_0_in [7]),
        .O(\r3/p_0_out [71]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[71]_i_1__2 
       (.I0(\r4/t0/t3/p_1_in [7]),
        .I1(\r4/t2/t1/p_0_in [7]),
        .I2(\r4/t1/t0/p_1_in [7]),
        .I3(\r4/t1/t0/p_0_in [7]),
        .I4(k3b[71]),
        .I5(\r4/t3/t2/p_0_in [7]),
        .O(\r4/p_0_out [71]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[71]_i_1__3 
       (.I0(\r5/t0/t3/p_1_in [7]),
        .I1(\r5/t2/t1/p_0_in [7]),
        .I2(\r5/t1/t0/p_1_in [7]),
        .I3(\r5/t1/t0/p_0_in [7]),
        .I4(k4b[71]),
        .I5(\r5/t3/t2/p_0_in [7]),
        .O(\r5/p_0_out [71]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[71]_i_1__4 
       (.I0(\r6/t0/t3/p_1_in [7]),
        .I1(\r6/t2/t1/p_0_in [7]),
        .I2(\r6/t1/t0/p_1_in [7]),
        .I3(\r6/t1/t0/p_0_in [7]),
        .I4(k5b[71]),
        .I5(\r6/t3/t2/p_0_in [7]),
        .O(\r6/p_0_out [71]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[71]_i_1__5 
       (.I0(\r7/t0/t3/p_1_in [7]),
        .I1(\r7/t2/t1/p_0_in [7]),
        .I2(\r7/t1/t0/p_1_in [7]),
        .I3(\r7/t1/t0/p_0_in [7]),
        .I4(k6b[71]),
        .I5(\r7/t3/t2/p_0_in [7]),
        .O(\r7/p_0_out [71]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[71]_i_1__6 
       (.I0(\r8/t0/t3/p_1_in [7]),
        .I1(\r8/t2/t1/p_0_in [7]),
        .I2(\r8/t1/t0/p_1_in [7]),
        .I3(\r8/t1/t0/p_0_in [7]),
        .I4(k7b[71]),
        .I5(\r8/t3/t2/p_0_in [7]),
        .O(\r8/p_0_out [71]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[71]_i_1__7 
       (.I0(\r9/t0/t3/p_1_in [7]),
        .I1(\r9/t2/t1/p_0_in [7]),
        .I2(\r9/t1/t0/p_1_in [7]),
        .I3(\r9/t1/t0/p_0_in [7]),
        .I4(k8b[71]),
        .I5(\r9/t3/t2/p_0_in [7]),
        .O(\r9/p_0_out [71]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair367" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[71]_i_1__8 
       (.I0(\a10/k1a [7]),
        .I1(\a10/k4a [7]),
        .I2(\rf/p_2_in [7]),
        .O(\rf/p_4_out [71]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[72]_i_1 
       (.I0(\r1/t0/t3/p_1_in [0]),
        .I1(\r1/t0/t3/p_0_in [0]),
        .I2(\r1/t2/t1/p_0_in [0]),
        .I3(\r1/t1/t0/p_0_in [0]),
        .I4(k0b[72]),
        .I5(\r1/t3/t2/p_1_in [0]),
        .O(\r1/p_0_out [72]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[72]_i_1__0 
       (.I0(\r2/t0/t3/p_1_in [0]),
        .I1(\r2/t0/t3/p_0_in [0]),
        .I2(\r2/t2/t1/p_0_in [0]),
        .I3(\r2/t1/t0/p_0_in [0]),
        .I4(k1b[72]),
        .I5(\r2/t3/t2/p_1_in [0]),
        .O(\r2/p_0_out [72]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[72]_i_1__1 
       (.I0(\r3/t0/t3/p_1_in [0]),
        .I1(\r3/t0/t3/p_0_in [0]),
        .I2(\r3/t2/t1/p_0_in [0]),
        .I3(\r3/t1/t0/p_0_in [0]),
        .I4(k2b[72]),
        .I5(\r3/t3/t2/p_1_in [0]),
        .O(\r3/p_0_out [72]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[72]_i_1__2 
       (.I0(\r4/t0/t3/p_1_in [0]),
        .I1(\r4/t0/t3/p_0_in [0]),
        .I2(\r4/t2/t1/p_0_in [0]),
        .I3(\r4/t1/t0/p_0_in [0]),
        .I4(k3b[72]),
        .I5(\r4/t3/t2/p_1_in [0]),
        .O(\r4/p_0_out [72]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[72]_i_1__3 
       (.I0(\r5/t0/t3/p_1_in [0]),
        .I1(\r5/t0/t3/p_0_in [0]),
        .I2(\r5/t2/t1/p_0_in [0]),
        .I3(\r5/t1/t0/p_0_in [0]),
        .I4(k4b[72]),
        .I5(\r5/t3/t2/p_1_in [0]),
        .O(\r5/p_0_out [72]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[72]_i_1__4 
       (.I0(\r6/t0/t3/p_1_in [0]),
        .I1(\r6/t0/t3/p_0_in [0]),
        .I2(\r6/t2/t1/p_0_in [0]),
        .I3(\r6/t1/t0/p_0_in [0]),
        .I4(k5b[72]),
        .I5(\r6/t3/t2/p_1_in [0]),
        .O(\r6/p_0_out [72]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[72]_i_1__5 
       (.I0(\r7/t0/t3/p_1_in [0]),
        .I1(\r7/t0/t3/p_0_in [0]),
        .I2(\r7/t2/t1/p_0_in [0]),
        .I3(\r7/t1/t0/p_0_in [0]),
        .I4(k6b[72]),
        .I5(\r7/t3/t2/p_1_in [0]),
        .O(\r7/p_0_out [72]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[72]_i_1__6 
       (.I0(\r8/t0/t3/p_1_in [0]),
        .I1(\r8/t0/t3/p_0_in [0]),
        .I2(\r8/t2/t1/p_0_in [0]),
        .I3(\r8/t1/t0/p_0_in [0]),
        .I4(k7b[72]),
        .I5(\r8/t3/t2/p_1_in [0]),
        .O(\r8/p_0_out [72]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[72]_i_1__7 
       (.I0(\r9/t0/t3/p_1_in [0]),
        .I1(\r9/t0/t3/p_0_in [0]),
        .I2(\r9/t2/t1/p_0_in [0]),
        .I3(\r9/t1/t0/p_0_in [0]),
        .I4(k8b[72]),
        .I5(\r9/t3/t2/p_1_in [0]),
        .O(\r9/p_0_out [72]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair366" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[72]_i_1__8 
       (.I0(\a10/k1a [8]),
        .I1(\a10/k4a [8]),
        .I2(\rf/p_2_in [8]),
        .O(\rf/p_4_out [72]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[73]_i_1 
       (.I0(\r1/t0/t3/p_1_in [1]),
        .I1(\r1/t0/t3/p_0_in [1]),
        .I2(\r1/t2/t1/p_0_in [1]),
        .I3(\r1/t1/t0/p_0_in [1]),
        .I4(k0b[73]),
        .I5(\r1/t3/t2/p_1_in [1]),
        .O(\r1/p_0_out [73]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[73]_i_1__0 
       (.I0(\r2/t0/t3/p_1_in [1]),
        .I1(\r2/t0/t3/p_0_in [1]),
        .I2(\r2/t2/t1/p_0_in [1]),
        .I3(\r2/t1/t0/p_0_in [1]),
        .I4(k1b[73]),
        .I5(\r2/t3/t2/p_1_in [1]),
        .O(\r2/p_0_out [73]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[73]_i_1__1 
       (.I0(\r3/t0/t3/p_1_in [1]),
        .I1(\r3/t0/t3/p_0_in [1]),
        .I2(\r3/t2/t1/p_0_in [1]),
        .I3(\r3/t1/t0/p_0_in [1]),
        .I4(k2b[73]),
        .I5(\r3/t3/t2/p_1_in [1]),
        .O(\r3/p_0_out [73]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[73]_i_1__2 
       (.I0(\r4/t0/t3/p_1_in [1]),
        .I1(\r4/t0/t3/p_0_in [1]),
        .I2(\r4/t2/t1/p_0_in [1]),
        .I3(\r4/t1/t0/p_0_in [1]),
        .I4(k3b[73]),
        .I5(\r4/t3/t2/p_1_in [1]),
        .O(\r4/p_0_out [73]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[73]_i_1__3 
       (.I0(\r5/t0/t3/p_1_in [1]),
        .I1(\r5/t0/t3/p_0_in [1]),
        .I2(\r5/t2/t1/p_0_in [1]),
        .I3(\r5/t1/t0/p_0_in [1]),
        .I4(k4b[73]),
        .I5(\r5/t3/t2/p_1_in [1]),
        .O(\r5/p_0_out [73]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[73]_i_1__4 
       (.I0(\r6/t0/t3/p_1_in [1]),
        .I1(\r6/t0/t3/p_0_in [1]),
        .I2(\r6/t2/t1/p_0_in [1]),
        .I3(\r6/t1/t0/p_0_in [1]),
        .I4(k5b[73]),
        .I5(\r6/t3/t2/p_1_in [1]),
        .O(\r6/p_0_out [73]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[73]_i_1__5 
       (.I0(\r7/t0/t3/p_1_in [1]),
        .I1(\r7/t0/t3/p_0_in [1]),
        .I2(\r7/t2/t1/p_0_in [1]),
        .I3(\r7/t1/t0/p_0_in [1]),
        .I4(k6b[73]),
        .I5(\r7/t3/t2/p_1_in [1]),
        .O(\r7/p_0_out [73]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[73]_i_1__6 
       (.I0(\r8/t0/t3/p_1_in [1]),
        .I1(\r8/t0/t3/p_0_in [1]),
        .I2(\r8/t2/t1/p_0_in [1]),
        .I3(\r8/t1/t0/p_0_in [1]),
        .I4(k7b[73]),
        .I5(\r8/t3/t2/p_1_in [1]),
        .O(\r8/p_0_out [73]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[73]_i_1__7 
       (.I0(\r9/t0/t3/p_1_in [1]),
        .I1(\r9/t0/t3/p_0_in [1]),
        .I2(\r9/t2/t1/p_0_in [1]),
        .I3(\r9/t1/t0/p_0_in [1]),
        .I4(k8b[73]),
        .I5(\r9/t3/t2/p_1_in [1]),
        .O(\r9/p_0_out [73]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair365" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[73]_i_1__8 
       (.I0(\a10/k1a [9]),
        .I1(\a10/k4a [9]),
        .I2(\rf/p_2_in [9]),
        .O(\rf/p_4_out [73]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[74]_i_1 
       (.I0(\r1/t0/t3/p_1_in [2]),
        .I1(\r1/t0/t3/p_0_in [2]),
        .I2(\r1/t2/t1/p_0_in [2]),
        .I3(\r1/t1/t0/p_0_in [2]),
        .I4(k0b[74]),
        .I5(\r1/t3/t2/p_1_in [2]),
        .O(\r1/p_0_out [74]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[74]_i_1__0 
       (.I0(\r2/t0/t3/p_1_in [2]),
        .I1(\r2/t0/t3/p_0_in [2]),
        .I2(\r2/t2/t1/p_0_in [2]),
        .I3(\r2/t1/t0/p_0_in [2]),
        .I4(k1b[74]),
        .I5(\r2/t3/t2/p_1_in [2]),
        .O(\r2/p_0_out [74]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[74]_i_1__1 
       (.I0(\r3/t0/t3/p_1_in [2]),
        .I1(\r3/t0/t3/p_0_in [2]),
        .I2(\r3/t2/t1/p_0_in [2]),
        .I3(\r3/t1/t0/p_0_in [2]),
        .I4(k2b[74]),
        .I5(\r3/t3/t2/p_1_in [2]),
        .O(\r3/p_0_out [74]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[74]_i_1__2 
       (.I0(\r4/t0/t3/p_1_in [2]),
        .I1(\r4/t0/t3/p_0_in [2]),
        .I2(\r4/t2/t1/p_0_in [2]),
        .I3(\r4/t1/t0/p_0_in [2]),
        .I4(k3b[74]),
        .I5(\r4/t3/t2/p_1_in [2]),
        .O(\r4/p_0_out [74]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[74]_i_1__3 
       (.I0(\r5/t0/t3/p_1_in [2]),
        .I1(\r5/t0/t3/p_0_in [2]),
        .I2(\r5/t2/t1/p_0_in [2]),
        .I3(\r5/t1/t0/p_0_in [2]),
        .I4(k4b[74]),
        .I5(\r5/t3/t2/p_1_in [2]),
        .O(\r5/p_0_out [74]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[74]_i_1__4 
       (.I0(\r6/t0/t3/p_1_in [2]),
        .I1(\r6/t0/t3/p_0_in [2]),
        .I2(\r6/t2/t1/p_0_in [2]),
        .I3(\r6/t1/t0/p_0_in [2]),
        .I4(k5b[74]),
        .I5(\r6/t3/t2/p_1_in [2]),
        .O(\r6/p_0_out [74]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[74]_i_1__5 
       (.I0(\r7/t0/t3/p_1_in [2]),
        .I1(\r7/t0/t3/p_0_in [2]),
        .I2(\r7/t2/t1/p_0_in [2]),
        .I3(\r7/t1/t0/p_0_in [2]),
        .I4(k6b[74]),
        .I5(\r7/t3/t2/p_1_in [2]),
        .O(\r7/p_0_out [74]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[74]_i_1__6 
       (.I0(\r8/t0/t3/p_1_in [2]),
        .I1(\r8/t0/t3/p_0_in [2]),
        .I2(\r8/t2/t1/p_0_in [2]),
        .I3(\r8/t1/t0/p_0_in [2]),
        .I4(k7b[74]),
        .I5(\r8/t3/t2/p_1_in [2]),
        .O(\r8/p_0_out [74]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[74]_i_1__7 
       (.I0(\r9/t0/t3/p_1_in [2]),
        .I1(\r9/t0/t3/p_0_in [2]),
        .I2(\r9/t2/t1/p_0_in [2]),
        .I3(\r9/t1/t0/p_0_in [2]),
        .I4(k8b[74]),
        .I5(\r9/t3/t2/p_1_in [2]),
        .O(\r9/p_0_out [74]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair364" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[74]_i_1__8 
       (.I0(\a10/k1a [10]),
        .I1(\a10/k4a [10]),
        .I2(\rf/p_2_in [10]),
        .O(\rf/p_4_out [74]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[75]_i_1 
       (.I0(\r1/t0/t3/p_1_in [3]),
        .I1(\r1/t0/t3/p_0_in [3]),
        .I2(\r1/t2/t1/p_0_in [3]),
        .I3(\r1/t1/t0/p_0_in [3]),
        .I4(k0b[75]),
        .I5(\r1/t3/t2/p_1_in [3]),
        .O(\r1/p_0_out [75]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[75]_i_1__0 
       (.I0(\r2/t0/t3/p_1_in [3]),
        .I1(\r2/t0/t3/p_0_in [3]),
        .I2(\r2/t2/t1/p_0_in [3]),
        .I3(\r2/t1/t0/p_0_in [3]),
        .I4(k1b[75]),
        .I5(\r2/t3/t2/p_1_in [3]),
        .O(\r2/p_0_out [75]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[75]_i_1__1 
       (.I0(\r3/t0/t3/p_1_in [3]),
        .I1(\r3/t0/t3/p_0_in [3]),
        .I2(\r3/t2/t1/p_0_in [3]),
        .I3(\r3/t1/t0/p_0_in [3]),
        .I4(k2b[75]),
        .I5(\r3/t3/t2/p_1_in [3]),
        .O(\r3/p_0_out [75]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[75]_i_1__2 
       (.I0(\r4/t0/t3/p_1_in [3]),
        .I1(\r4/t0/t3/p_0_in [3]),
        .I2(\r4/t2/t1/p_0_in [3]),
        .I3(\r4/t1/t0/p_0_in [3]),
        .I4(k3b[75]),
        .I5(\r4/t3/t2/p_1_in [3]),
        .O(\r4/p_0_out [75]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[75]_i_1__3 
       (.I0(\r5/t0/t3/p_1_in [3]),
        .I1(\r5/t0/t3/p_0_in [3]),
        .I2(\r5/t2/t1/p_0_in [3]),
        .I3(\r5/t1/t0/p_0_in [3]),
        .I4(k4b[75]),
        .I5(\r5/t3/t2/p_1_in [3]),
        .O(\r5/p_0_out [75]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[75]_i_1__4 
       (.I0(\r6/t0/t3/p_1_in [3]),
        .I1(\r6/t0/t3/p_0_in [3]),
        .I2(\r6/t2/t1/p_0_in [3]),
        .I3(\r6/t1/t0/p_0_in [3]),
        .I4(k5b[75]),
        .I5(\r6/t3/t2/p_1_in [3]),
        .O(\r6/p_0_out [75]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[75]_i_1__5 
       (.I0(\r7/t0/t3/p_1_in [3]),
        .I1(\r7/t0/t3/p_0_in [3]),
        .I2(\r7/t2/t1/p_0_in [3]),
        .I3(\r7/t1/t0/p_0_in [3]),
        .I4(k6b[75]),
        .I5(\r7/t3/t2/p_1_in [3]),
        .O(\r7/p_0_out [75]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[75]_i_1__6 
       (.I0(\r8/t0/t3/p_1_in [3]),
        .I1(\r8/t0/t3/p_0_in [3]),
        .I2(\r8/t2/t1/p_0_in [3]),
        .I3(\r8/t1/t0/p_0_in [3]),
        .I4(k7b[75]),
        .I5(\r8/t3/t2/p_1_in [3]),
        .O(\r8/p_0_out [75]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[75]_i_1__7 
       (.I0(\r9/t0/t3/p_1_in [3]),
        .I1(\r9/t0/t3/p_0_in [3]),
        .I2(\r9/t2/t1/p_0_in [3]),
        .I3(\r9/t1/t0/p_0_in [3]),
        .I4(k8b[75]),
        .I5(\r9/t3/t2/p_1_in [3]),
        .O(\r9/p_0_out [75]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair363" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[75]_i_1__8 
       (.I0(\a10/k1a [11]),
        .I1(\a10/k4a [11]),
        .I2(\rf/p_2_in [11]),
        .O(\rf/p_4_out [75]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[76]_i_1 
       (.I0(\r1/t0/t3/p_1_in [4]),
        .I1(\r1/t0/t3/p_0_in [4]),
        .I2(\r1/t2/t1/p_0_in [4]),
        .I3(\r1/t1/t0/p_0_in [4]),
        .I4(k0b[76]),
        .I5(\r1/t3/t2/p_1_in [4]),
        .O(\r1/p_0_out [76]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[76]_i_1__0 
       (.I0(\r2/t0/t3/p_1_in [4]),
        .I1(\r2/t0/t3/p_0_in [4]),
        .I2(\r2/t2/t1/p_0_in [4]),
        .I3(\r2/t1/t0/p_0_in [4]),
        .I4(k1b[76]),
        .I5(\r2/t3/t2/p_1_in [4]),
        .O(\r2/p_0_out [76]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[76]_i_1__1 
       (.I0(\r3/t0/t3/p_1_in [4]),
        .I1(\r3/t0/t3/p_0_in [4]),
        .I2(\r3/t2/t1/p_0_in [4]),
        .I3(\r3/t1/t0/p_0_in [4]),
        .I4(k2b[76]),
        .I5(\r3/t3/t2/p_1_in [4]),
        .O(\r3/p_0_out [76]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[76]_i_1__2 
       (.I0(\r4/t0/t3/p_1_in [4]),
        .I1(\r4/t0/t3/p_0_in [4]),
        .I2(\r4/t2/t1/p_0_in [4]),
        .I3(\r4/t1/t0/p_0_in [4]),
        .I4(k3b[76]),
        .I5(\r4/t3/t2/p_1_in [4]),
        .O(\r4/p_0_out [76]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[76]_i_1__3 
       (.I0(\r5/t0/t3/p_1_in [4]),
        .I1(\r5/t0/t3/p_0_in [4]),
        .I2(\r5/t2/t1/p_0_in [4]),
        .I3(\r5/t1/t0/p_0_in [4]),
        .I4(k4b[76]),
        .I5(\r5/t3/t2/p_1_in [4]),
        .O(\r5/p_0_out [76]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[76]_i_1__4 
       (.I0(\r6/t0/t3/p_1_in [4]),
        .I1(\r6/t0/t3/p_0_in [4]),
        .I2(\r6/t2/t1/p_0_in [4]),
        .I3(\r6/t1/t0/p_0_in [4]),
        .I4(k5b[76]),
        .I5(\r6/t3/t2/p_1_in [4]),
        .O(\r6/p_0_out [76]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[76]_i_1__5 
       (.I0(\r7/t0/t3/p_1_in [4]),
        .I1(\r7/t0/t3/p_0_in [4]),
        .I2(\r7/t2/t1/p_0_in [4]),
        .I3(\r7/t1/t0/p_0_in [4]),
        .I4(k6b[76]),
        .I5(\r7/t3/t2/p_1_in [4]),
        .O(\r7/p_0_out [76]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[76]_i_1__6 
       (.I0(\r8/t0/t3/p_1_in [4]),
        .I1(\r8/t0/t3/p_0_in [4]),
        .I2(\r8/t2/t1/p_0_in [4]),
        .I3(\r8/t1/t0/p_0_in [4]),
        .I4(k7b[76]),
        .I5(\r8/t3/t2/p_1_in [4]),
        .O(\r8/p_0_out [76]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[76]_i_1__7 
       (.I0(\r9/t0/t3/p_1_in [4]),
        .I1(\r9/t0/t3/p_0_in [4]),
        .I2(\r9/t2/t1/p_0_in [4]),
        .I3(\r9/t1/t0/p_0_in [4]),
        .I4(k8b[76]),
        .I5(\r9/t3/t2/p_1_in [4]),
        .O(\r9/p_0_out [76]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair362" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[76]_i_1__8 
       (.I0(\a10/k1a [12]),
        .I1(\a10/k4a [12]),
        .I2(\rf/p_2_in [12]),
        .O(\rf/p_4_out [76]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[77]_i_1 
       (.I0(\r1/t0/t3/p_1_in [5]),
        .I1(\r1/t0/t3/p_0_in [5]),
        .I2(\r1/t2/t1/p_0_in [5]),
        .I3(\r1/t1/t0/p_0_in [5]),
        .I4(k0b[77]),
        .I5(\r1/t3/t2/p_1_in [5]),
        .O(\r1/p_0_out [77]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[77]_i_1__0 
       (.I0(\r2/t0/t3/p_1_in [5]),
        .I1(\r2/t0/t3/p_0_in [5]),
        .I2(\r2/t2/t1/p_0_in [5]),
        .I3(\r2/t1/t0/p_0_in [5]),
        .I4(k1b[77]),
        .I5(\r2/t3/t2/p_1_in [5]),
        .O(\r2/p_0_out [77]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[77]_i_1__1 
       (.I0(\r3/t0/t3/p_1_in [5]),
        .I1(\r3/t0/t3/p_0_in [5]),
        .I2(\r3/t2/t1/p_0_in [5]),
        .I3(\r3/t1/t0/p_0_in [5]),
        .I4(k2b[77]),
        .I5(\r3/t3/t2/p_1_in [5]),
        .O(\r3/p_0_out [77]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[77]_i_1__2 
       (.I0(\r4/t0/t3/p_1_in [5]),
        .I1(\r4/t0/t3/p_0_in [5]),
        .I2(\r4/t2/t1/p_0_in [5]),
        .I3(\r4/t1/t0/p_0_in [5]),
        .I4(k3b[77]),
        .I5(\r4/t3/t2/p_1_in [5]),
        .O(\r4/p_0_out [77]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[77]_i_1__3 
       (.I0(\r5/t0/t3/p_1_in [5]),
        .I1(\r5/t0/t3/p_0_in [5]),
        .I2(\r5/t2/t1/p_0_in [5]),
        .I3(\r5/t1/t0/p_0_in [5]),
        .I4(k4b[77]),
        .I5(\r5/t3/t2/p_1_in [5]),
        .O(\r5/p_0_out [77]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[77]_i_1__4 
       (.I0(\r6/t0/t3/p_1_in [5]),
        .I1(\r6/t0/t3/p_0_in [5]),
        .I2(\r6/t2/t1/p_0_in [5]),
        .I3(\r6/t1/t0/p_0_in [5]),
        .I4(k5b[77]),
        .I5(\r6/t3/t2/p_1_in [5]),
        .O(\r6/p_0_out [77]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[77]_i_1__5 
       (.I0(\r7/t0/t3/p_1_in [5]),
        .I1(\r7/t0/t3/p_0_in [5]),
        .I2(\r7/t2/t1/p_0_in [5]),
        .I3(\r7/t1/t0/p_0_in [5]),
        .I4(k6b[77]),
        .I5(\r7/t3/t2/p_1_in [5]),
        .O(\r7/p_0_out [77]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[77]_i_1__6 
       (.I0(\r8/t0/t3/p_1_in [5]),
        .I1(\r8/t0/t3/p_0_in [5]),
        .I2(\r8/t2/t1/p_0_in [5]),
        .I3(\r8/t1/t0/p_0_in [5]),
        .I4(k7b[77]),
        .I5(\r8/t3/t2/p_1_in [5]),
        .O(\r8/p_0_out [77]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[77]_i_1__7 
       (.I0(\r9/t0/t3/p_1_in [5]),
        .I1(\r9/t0/t3/p_0_in [5]),
        .I2(\r9/t2/t1/p_0_in [5]),
        .I3(\r9/t1/t0/p_0_in [5]),
        .I4(k8b[77]),
        .I5(\r9/t3/t2/p_1_in [5]),
        .O(\r9/p_0_out [77]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair361" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[77]_i_1__8 
       (.I0(\a10/k1a [13]),
        .I1(\a10/k4a [13]),
        .I2(\rf/p_2_in [13]),
        .O(\rf/p_4_out [77]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[78]_i_1 
       (.I0(\r1/t0/t3/p_1_in [6]),
        .I1(\r1/t0/t3/p_0_in [6]),
        .I2(\r1/t2/t1/p_0_in [6]),
        .I3(\r1/t1/t0/p_0_in [6]),
        .I4(k0b[78]),
        .I5(\r1/t3/t2/p_1_in [6]),
        .O(\r1/p_0_out [78]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[78]_i_1__0 
       (.I0(\r2/t0/t3/p_1_in [6]),
        .I1(\r2/t0/t3/p_0_in [6]),
        .I2(\r2/t2/t1/p_0_in [6]),
        .I3(\r2/t1/t0/p_0_in [6]),
        .I4(k1b[78]),
        .I5(\r2/t3/t2/p_1_in [6]),
        .O(\r2/p_0_out [78]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[78]_i_1__1 
       (.I0(\r3/t0/t3/p_1_in [6]),
        .I1(\r3/t0/t3/p_0_in [6]),
        .I2(\r3/t2/t1/p_0_in [6]),
        .I3(\r3/t1/t0/p_0_in [6]),
        .I4(k2b[78]),
        .I5(\r3/t3/t2/p_1_in [6]),
        .O(\r3/p_0_out [78]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[78]_i_1__2 
       (.I0(\r4/t0/t3/p_1_in [6]),
        .I1(\r4/t0/t3/p_0_in [6]),
        .I2(\r4/t2/t1/p_0_in [6]),
        .I3(\r4/t1/t0/p_0_in [6]),
        .I4(k3b[78]),
        .I5(\r4/t3/t2/p_1_in [6]),
        .O(\r4/p_0_out [78]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[78]_i_1__3 
       (.I0(\r5/t0/t3/p_1_in [6]),
        .I1(\r5/t0/t3/p_0_in [6]),
        .I2(\r5/t2/t1/p_0_in [6]),
        .I3(\r5/t1/t0/p_0_in [6]),
        .I4(k4b[78]),
        .I5(\r5/t3/t2/p_1_in [6]),
        .O(\r5/p_0_out [78]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[78]_i_1__4 
       (.I0(\r6/t0/t3/p_1_in [6]),
        .I1(\r6/t0/t3/p_0_in [6]),
        .I2(\r6/t2/t1/p_0_in [6]),
        .I3(\r6/t1/t0/p_0_in [6]),
        .I4(k5b[78]),
        .I5(\r6/t3/t2/p_1_in [6]),
        .O(\r6/p_0_out [78]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[78]_i_1__5 
       (.I0(\r7/t0/t3/p_1_in [6]),
        .I1(\r7/t0/t3/p_0_in [6]),
        .I2(\r7/t2/t1/p_0_in [6]),
        .I3(\r7/t1/t0/p_0_in [6]),
        .I4(k6b[78]),
        .I5(\r7/t3/t2/p_1_in [6]),
        .O(\r7/p_0_out [78]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[78]_i_1__6 
       (.I0(\r8/t0/t3/p_1_in [6]),
        .I1(\r8/t0/t3/p_0_in [6]),
        .I2(\r8/t2/t1/p_0_in [6]),
        .I3(\r8/t1/t0/p_0_in [6]),
        .I4(k7b[78]),
        .I5(\r8/t3/t2/p_1_in [6]),
        .O(\r8/p_0_out [78]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[78]_i_1__7 
       (.I0(\r9/t0/t3/p_1_in [6]),
        .I1(\r9/t0/t3/p_0_in [6]),
        .I2(\r9/t2/t1/p_0_in [6]),
        .I3(\r9/t1/t0/p_0_in [6]),
        .I4(k8b[78]),
        .I5(\r9/t3/t2/p_1_in [6]),
        .O(\r9/p_0_out [78]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair383" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[78]_i_1__8 
       (.I0(\a10/k1a [14]),
        .I1(\a10/k4a [14]),
        .I2(\rf/p_2_in [14]),
        .O(\rf/p_4_out [78]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[79]_i_1 
       (.I0(\r1/t0/t3/p_1_in [7]),
        .I1(\r1/t0/t3/p_0_in [7]),
        .I2(\r1/t2/t1/p_0_in [7]),
        .I3(\r1/t1/t0/p_0_in [7]),
        .I4(k0b[79]),
        .I5(\r1/t3/t2/p_1_in [7]),
        .O(\r1/p_0_out [79]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[79]_i_1__0 
       (.I0(\r2/t0/t3/p_1_in [7]),
        .I1(\r2/t0/t3/p_0_in [7]),
        .I2(\r2/t2/t1/p_0_in [7]),
        .I3(\r2/t1/t0/p_0_in [7]),
        .I4(k1b[79]),
        .I5(\r2/t3/t2/p_1_in [7]),
        .O(\r2/p_0_out [79]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[79]_i_1__1 
       (.I0(\r3/t0/t3/p_1_in [7]),
        .I1(\r3/t0/t3/p_0_in [7]),
        .I2(\r3/t2/t1/p_0_in [7]),
        .I3(\r3/t1/t0/p_0_in [7]),
        .I4(k2b[79]),
        .I5(\r3/t3/t2/p_1_in [7]),
        .O(\r3/p_0_out [79]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[79]_i_1__2 
       (.I0(\r4/t0/t3/p_1_in [7]),
        .I1(\r4/t0/t3/p_0_in [7]),
        .I2(\r4/t2/t1/p_0_in [7]),
        .I3(\r4/t1/t0/p_0_in [7]),
        .I4(k3b[79]),
        .I5(\r4/t3/t2/p_1_in [7]),
        .O(\r4/p_0_out [79]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[79]_i_1__3 
       (.I0(\r5/t0/t3/p_1_in [7]),
        .I1(\r5/t0/t3/p_0_in [7]),
        .I2(\r5/t2/t1/p_0_in [7]),
        .I3(\r5/t1/t0/p_0_in [7]),
        .I4(k4b[79]),
        .I5(\r5/t3/t2/p_1_in [7]),
        .O(\r5/p_0_out [79]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[79]_i_1__4 
       (.I0(\r6/t0/t3/p_1_in [7]),
        .I1(\r6/t0/t3/p_0_in [7]),
        .I2(\r6/t2/t1/p_0_in [7]),
        .I3(\r6/t1/t0/p_0_in [7]),
        .I4(k5b[79]),
        .I5(\r6/t3/t2/p_1_in [7]),
        .O(\r6/p_0_out [79]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[79]_i_1__5 
       (.I0(\r7/t0/t3/p_1_in [7]),
        .I1(\r7/t0/t3/p_0_in [7]),
        .I2(\r7/t2/t1/p_0_in [7]),
        .I3(\r7/t1/t0/p_0_in [7]),
        .I4(k6b[79]),
        .I5(\r7/t3/t2/p_1_in [7]),
        .O(\r7/p_0_out [79]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[79]_i_1__6 
       (.I0(\r8/t0/t3/p_1_in [7]),
        .I1(\r8/t0/t3/p_0_in [7]),
        .I2(\r8/t2/t1/p_0_in [7]),
        .I3(\r8/t1/t0/p_0_in [7]),
        .I4(k7b[79]),
        .I5(\r8/t3/t2/p_1_in [7]),
        .O(\r8/p_0_out [79]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[79]_i_1__7 
       (.I0(\r9/t0/t3/p_1_in [7]),
        .I1(\r9/t0/t3/p_0_in [7]),
        .I2(\r9/t2/t1/p_0_in [7]),
        .I3(\r9/t1/t0/p_0_in [7]),
        .I4(k8b[79]),
        .I5(\r9/t3/t2/p_1_in [7]),
        .O(\r9/p_0_out [79]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair359" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[79]_i_1__8 
       (.I0(\a10/k1a [15]),
        .I1(\a10/k4a [15]),
        .I2(\rf/p_2_in [15]),
        .O(\rf/p_4_out [79]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[7]_i_1 
       (.I0(\r1/t0/t1/p_0_in [7]),
        .I1(\r1/t2/t3/p_1_in [7]),
        .I2(\r1/t1/t2/p_0_in [7]),
        .I3(k0b[7]),
        .I4(\r1/t3/t0/p_1_in [7]),
        .I5(\r1/t3/t0/p_0_in [7]),
        .O(\r1/p_0_out [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[7]_i_1__0 
       (.I0(\r2/t0/t1/p_0_in [7]),
        .I1(\r2/t2/t3/p_1_in [7]),
        .I2(\r2/t1/t2/p_0_in [7]),
        .I3(k1b[7]),
        .I4(\r2/t3/t0/p_1_in [7]),
        .I5(\r2/t3/t0/p_0_in [7]),
        .O(\r2/p_0_out [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[7]_i_1__1 
       (.I0(\r3/t0/t1/p_0_in [7]),
        .I1(\r3/t2/t3/p_1_in [7]),
        .I2(\r3/t1/t2/p_0_in [7]),
        .I3(k2b[7]),
        .I4(\r3/t3/t0/p_1_in [7]),
        .I5(\r3/t3/t0/p_0_in [7]),
        .O(\r3/p_0_out [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[7]_i_1__2 
       (.I0(\r4/t0/t1/p_0_in [7]),
        .I1(\r4/t2/t3/p_1_in [7]),
        .I2(\r4/t1/t2/p_0_in [7]),
        .I3(k3b[7]),
        .I4(\r4/t3/t0/p_1_in [7]),
        .I5(\r4/t3/t0/p_0_in [7]),
        .O(\r4/p_0_out [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[7]_i_1__3 
       (.I0(\r5/t0/t1/p_0_in [7]),
        .I1(\r5/t2/t3/p_1_in [7]),
        .I2(\r5/t1/t2/p_0_in [7]),
        .I3(k4b[7]),
        .I4(\r5/t3/t0/p_1_in [7]),
        .I5(\r5/t3/t0/p_0_in [7]),
        .O(\r5/p_0_out [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[7]_i_1__4 
       (.I0(\r6/t0/t1/p_0_in [7]),
        .I1(\r6/t2/t3/p_1_in [7]),
        .I2(\r6/t1/t2/p_0_in [7]),
        .I3(k5b[7]),
        .I4(\r6/t3/t0/p_1_in [7]),
        .I5(\r6/t3/t0/p_0_in [7]),
        .O(\r6/p_0_out [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[7]_i_1__5 
       (.I0(\r7/t0/t1/p_0_in [7]),
        .I1(\r7/t2/t3/p_1_in [7]),
        .I2(\r7/t1/t2/p_0_in [7]),
        .I3(k6b[7]),
        .I4(\r7/t3/t0/p_1_in [7]),
        .I5(\r7/t3/t0/p_0_in [7]),
        .O(\r7/p_0_out [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[7]_i_1__6 
       (.I0(\r8/t0/t1/p_0_in [7]),
        .I1(\r8/t2/t3/p_1_in [7]),
        .I2(\r8/t1/t2/p_0_in [7]),
        .I3(k7b[7]),
        .I4(\r8/t3/t0/p_1_in [7]),
        .I5(\r8/t3/t0/p_0_in [7]),
        .O(\r8/p_0_out [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[7]_i_1__7 
       (.I0(\r9/t0/t1/p_0_in [7]),
        .I1(\r9/t2/t3/p_1_in [7]),
        .I2(\r9/t1/t2/p_0_in [7]),
        .I3(k8b[7]),
        .I4(\r9/t3/t0/p_1_in [7]),
        .I5(\r9/t3/t0/p_0_in [7]),
        .O(\r9/p_0_out [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair335" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[7]_i_1__8 
       (.I0(\a10/k3a [7]),
        .I1(\a10/k4a [7]),
        .I2(\rf/p_0_in [7]),
        .O(\rf/p_4_out [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[80]_i_1 
       (.I0(\r1/t0/t3/p_0_in [0]),
        .I1(\r1/t2/t1/p_1_in [0]),
        .I2(\r1/t1/t0/p_0_in [0]),
        .I3(k0b[80]),
        .I4(\r1/t3/t2/p_1_in [0]),
        .I5(\r1/t3/t2/p_0_in [0]),
        .O(\r1/p_0_out [80]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[80]_i_1__0 
       (.I0(\r2/t0/t3/p_0_in [0]),
        .I1(\r2/t2/t1/p_1_in [0]),
        .I2(\r2/t1/t0/p_0_in [0]),
        .I3(k1b[80]),
        .I4(\r2/t3/t2/p_1_in [0]),
        .I5(\r2/t3/t2/p_0_in [0]),
        .O(\r2/p_0_out [80]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[80]_i_1__1 
       (.I0(\r3/t0/t3/p_0_in [0]),
        .I1(\r3/t2/t1/p_1_in [0]),
        .I2(\r3/t1/t0/p_0_in [0]),
        .I3(k2b[80]),
        .I4(\r3/t3/t2/p_1_in [0]),
        .I5(\r3/t3/t2/p_0_in [0]),
        .O(\r3/p_0_out [80]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[80]_i_1__2 
       (.I0(\r4/t0/t3/p_0_in [0]),
        .I1(\r4/t2/t1/p_1_in [0]),
        .I2(\r4/t1/t0/p_0_in [0]),
        .I3(k3b[80]),
        .I4(\r4/t3/t2/p_1_in [0]),
        .I5(\r4/t3/t2/p_0_in [0]),
        .O(\r4/p_0_out [80]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[80]_i_1__3 
       (.I0(\r5/t0/t3/p_0_in [0]),
        .I1(\r5/t2/t1/p_1_in [0]),
        .I2(\r5/t1/t0/p_0_in [0]),
        .I3(k4b[80]),
        .I4(\r5/t3/t2/p_1_in [0]),
        .I5(\r5/t3/t2/p_0_in [0]),
        .O(\r5/p_0_out [80]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[80]_i_1__4 
       (.I0(\r6/t0/t3/p_0_in [0]),
        .I1(\r6/t2/t1/p_1_in [0]),
        .I2(\r6/t1/t0/p_0_in [0]),
        .I3(k5b[80]),
        .I4(\r6/t3/t2/p_1_in [0]),
        .I5(\r6/t3/t2/p_0_in [0]),
        .O(\r6/p_0_out [80]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[80]_i_1__5 
       (.I0(\r7/t0/t3/p_0_in [0]),
        .I1(\r7/t2/t1/p_1_in [0]),
        .I2(\r7/t1/t0/p_0_in [0]),
        .I3(k6b[80]),
        .I4(\r7/t3/t2/p_1_in [0]),
        .I5(\r7/t3/t2/p_0_in [0]),
        .O(\r7/p_0_out [80]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[80]_i_1__6 
       (.I0(\r8/t0/t3/p_0_in [0]),
        .I1(\r8/t2/t1/p_1_in [0]),
        .I2(\r8/t1/t0/p_0_in [0]),
        .I3(k7b[80]),
        .I4(\r8/t3/t2/p_1_in [0]),
        .I5(\r8/t3/t2/p_0_in [0]),
        .O(\r8/p_0_out [80]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[80]_i_1__7 
       (.I0(\r9/t0/t3/p_0_in [0]),
        .I1(\r9/t2/t1/p_1_in [0]),
        .I2(\r9/t1/t0/p_0_in [0]),
        .I3(k8b[80]),
        .I4(\r9/t3/t2/p_1_in [0]),
        .I5(\r9/t3/t2/p_0_in [0]),
        .O(\r9/p_0_out [80]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair358" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[80]_i_1__8 
       (.I0(\a10/k1a [16]),
        .I1(\a10/k4a [16]),
        .I2(\rf/p_2_in [16]),
        .O(\rf/p_4_out [80]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[81]_i_1 
       (.I0(\r1/t0/t3/p_0_in [1]),
        .I1(\r1/t2/t1/p_1_in [1]),
        .I2(\r1/t1/t0/p_0_in [1]),
        .I3(k0b[81]),
        .I4(\r1/t3/t2/p_1_in [1]),
        .I5(\r1/t3/t2/p_0_in [1]),
        .O(\r1/p_0_out [81]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[81]_i_1__0 
       (.I0(\r2/t0/t3/p_0_in [1]),
        .I1(\r2/t2/t1/p_1_in [1]),
        .I2(\r2/t1/t0/p_0_in [1]),
        .I3(k1b[81]),
        .I4(\r2/t3/t2/p_1_in [1]),
        .I5(\r2/t3/t2/p_0_in [1]),
        .O(\r2/p_0_out [81]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[81]_i_1__1 
       (.I0(\r3/t0/t3/p_0_in [1]),
        .I1(\r3/t2/t1/p_1_in [1]),
        .I2(\r3/t1/t0/p_0_in [1]),
        .I3(k2b[81]),
        .I4(\r3/t3/t2/p_1_in [1]),
        .I5(\r3/t3/t2/p_0_in [1]),
        .O(\r3/p_0_out [81]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[81]_i_1__2 
       (.I0(\r4/t0/t3/p_0_in [1]),
        .I1(\r4/t2/t1/p_1_in [1]),
        .I2(\r4/t1/t0/p_0_in [1]),
        .I3(k3b[81]),
        .I4(\r4/t3/t2/p_1_in [1]),
        .I5(\r4/t3/t2/p_0_in [1]),
        .O(\r4/p_0_out [81]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[81]_i_1__3 
       (.I0(\r5/t0/t3/p_0_in [1]),
        .I1(\r5/t2/t1/p_1_in [1]),
        .I2(\r5/t1/t0/p_0_in [1]),
        .I3(k4b[81]),
        .I4(\r5/t3/t2/p_1_in [1]),
        .I5(\r5/t3/t2/p_0_in [1]),
        .O(\r5/p_0_out [81]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[81]_i_1__4 
       (.I0(\r6/t0/t3/p_0_in [1]),
        .I1(\r6/t2/t1/p_1_in [1]),
        .I2(\r6/t1/t0/p_0_in [1]),
        .I3(k5b[81]),
        .I4(\r6/t3/t2/p_1_in [1]),
        .I5(\r6/t3/t2/p_0_in [1]),
        .O(\r6/p_0_out [81]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[81]_i_1__5 
       (.I0(\r7/t0/t3/p_0_in [1]),
        .I1(\r7/t2/t1/p_1_in [1]),
        .I2(\r7/t1/t0/p_0_in [1]),
        .I3(k6b[81]),
        .I4(\r7/t3/t2/p_1_in [1]),
        .I5(\r7/t3/t2/p_0_in [1]),
        .O(\r7/p_0_out [81]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[81]_i_1__6 
       (.I0(\r8/t0/t3/p_0_in [1]),
        .I1(\r8/t2/t1/p_1_in [1]),
        .I2(\r8/t1/t0/p_0_in [1]),
        .I3(k7b[81]),
        .I4(\r8/t3/t2/p_1_in [1]),
        .I5(\r8/t3/t2/p_0_in [1]),
        .O(\r8/p_0_out [81]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[81]_i_1__7 
       (.I0(\r9/t0/t3/p_0_in [1]),
        .I1(\r9/t2/t1/p_1_in [1]),
        .I2(\r9/t1/t0/p_0_in [1]),
        .I3(k8b[81]),
        .I4(\r9/t3/t2/p_1_in [1]),
        .I5(\r9/t3/t2/p_0_in [1]),
        .O(\r9/p_0_out [81]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair357" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[81]_i_1__8 
       (.I0(\a10/k1a [17]),
        .I1(\a10/k4a [17]),
        .I2(\rf/p_2_in [17]),
        .O(\rf/p_4_out [81]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[82]_i_1 
       (.I0(\r1/t0/t3/p_0_in [2]),
        .I1(\r1/t2/t1/p_1_in [2]),
        .I2(\r1/t1/t0/p_0_in [2]),
        .I3(k0b[82]),
        .I4(\r1/t3/t2/p_1_in [2]),
        .I5(\r1/t3/t2/p_0_in [2]),
        .O(\r1/p_0_out [82]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[82]_i_1__0 
       (.I0(\r2/t0/t3/p_0_in [2]),
        .I1(\r2/t2/t1/p_1_in [2]),
        .I2(\r2/t1/t0/p_0_in [2]),
        .I3(k1b[82]),
        .I4(\r2/t3/t2/p_1_in [2]),
        .I5(\r2/t3/t2/p_0_in [2]),
        .O(\r2/p_0_out [82]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[82]_i_1__1 
       (.I0(\r3/t0/t3/p_0_in [2]),
        .I1(\r3/t2/t1/p_1_in [2]),
        .I2(\r3/t1/t0/p_0_in [2]),
        .I3(k2b[82]),
        .I4(\r3/t3/t2/p_1_in [2]),
        .I5(\r3/t3/t2/p_0_in [2]),
        .O(\r3/p_0_out [82]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[82]_i_1__2 
       (.I0(\r4/t0/t3/p_0_in [2]),
        .I1(\r4/t2/t1/p_1_in [2]),
        .I2(\r4/t1/t0/p_0_in [2]),
        .I3(k3b[82]),
        .I4(\r4/t3/t2/p_1_in [2]),
        .I5(\r4/t3/t2/p_0_in [2]),
        .O(\r4/p_0_out [82]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[82]_i_1__3 
       (.I0(\r5/t0/t3/p_0_in [2]),
        .I1(\r5/t2/t1/p_1_in [2]),
        .I2(\r5/t1/t0/p_0_in [2]),
        .I3(k4b[82]),
        .I4(\r5/t3/t2/p_1_in [2]),
        .I5(\r5/t3/t2/p_0_in [2]),
        .O(\r5/p_0_out [82]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[82]_i_1__4 
       (.I0(\r6/t0/t3/p_0_in [2]),
        .I1(\r6/t2/t1/p_1_in [2]),
        .I2(\r6/t1/t0/p_0_in [2]),
        .I3(k5b[82]),
        .I4(\r6/t3/t2/p_1_in [2]),
        .I5(\r6/t3/t2/p_0_in [2]),
        .O(\r6/p_0_out [82]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[82]_i_1__5 
       (.I0(\r7/t0/t3/p_0_in [2]),
        .I1(\r7/t2/t1/p_1_in [2]),
        .I2(\r7/t1/t0/p_0_in [2]),
        .I3(k6b[82]),
        .I4(\r7/t3/t2/p_1_in [2]),
        .I5(\r7/t3/t2/p_0_in [2]),
        .O(\r7/p_0_out [82]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[82]_i_1__6 
       (.I0(\r8/t0/t3/p_0_in [2]),
        .I1(\r8/t2/t1/p_1_in [2]),
        .I2(\r8/t1/t0/p_0_in [2]),
        .I3(k7b[82]),
        .I4(\r8/t3/t2/p_1_in [2]),
        .I5(\r8/t3/t2/p_0_in [2]),
        .O(\r8/p_0_out [82]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[82]_i_1__7 
       (.I0(\r9/t0/t3/p_0_in [2]),
        .I1(\r9/t2/t1/p_1_in [2]),
        .I2(\r9/t1/t0/p_0_in [2]),
        .I3(k8b[82]),
        .I4(\r9/t3/t2/p_1_in [2]),
        .I5(\r9/t3/t2/p_0_in [2]),
        .O(\r9/p_0_out [82]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair356" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[82]_i_1__8 
       (.I0(\a10/k1a [18]),
        .I1(\a10/k4a [18]),
        .I2(\rf/p_2_in [18]),
        .O(\rf/p_4_out [82]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[83]_i_1 
       (.I0(\r1/t0/t3/p_0_in [3]),
        .I1(\r1/t2/t1/p_1_in [3]),
        .I2(\r1/t1/t0/p_0_in [3]),
        .I3(k0b[83]),
        .I4(\r1/t3/t2/p_1_in [3]),
        .I5(\r1/t3/t2/p_0_in [3]),
        .O(\r1/p_0_out [83]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[83]_i_1__0 
       (.I0(\r2/t0/t3/p_0_in [3]),
        .I1(\r2/t2/t1/p_1_in [3]),
        .I2(\r2/t1/t0/p_0_in [3]),
        .I3(k1b[83]),
        .I4(\r2/t3/t2/p_1_in [3]),
        .I5(\r2/t3/t2/p_0_in [3]),
        .O(\r2/p_0_out [83]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[83]_i_1__1 
       (.I0(\r3/t0/t3/p_0_in [3]),
        .I1(\r3/t2/t1/p_1_in [3]),
        .I2(\r3/t1/t0/p_0_in [3]),
        .I3(k2b[83]),
        .I4(\r3/t3/t2/p_1_in [3]),
        .I5(\r3/t3/t2/p_0_in [3]),
        .O(\r3/p_0_out [83]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[83]_i_1__2 
       (.I0(\r4/t0/t3/p_0_in [3]),
        .I1(\r4/t2/t1/p_1_in [3]),
        .I2(\r4/t1/t0/p_0_in [3]),
        .I3(k3b[83]),
        .I4(\r4/t3/t2/p_1_in [3]),
        .I5(\r4/t3/t2/p_0_in [3]),
        .O(\r4/p_0_out [83]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[83]_i_1__3 
       (.I0(\r5/t0/t3/p_0_in [3]),
        .I1(\r5/t2/t1/p_1_in [3]),
        .I2(\r5/t1/t0/p_0_in [3]),
        .I3(k4b[83]),
        .I4(\r5/t3/t2/p_1_in [3]),
        .I5(\r5/t3/t2/p_0_in [3]),
        .O(\r5/p_0_out [83]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[83]_i_1__4 
       (.I0(\r6/t0/t3/p_0_in [3]),
        .I1(\r6/t2/t1/p_1_in [3]),
        .I2(\r6/t1/t0/p_0_in [3]),
        .I3(k5b[83]),
        .I4(\r6/t3/t2/p_1_in [3]),
        .I5(\r6/t3/t2/p_0_in [3]),
        .O(\r6/p_0_out [83]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[83]_i_1__5 
       (.I0(\r7/t0/t3/p_0_in [3]),
        .I1(\r7/t2/t1/p_1_in [3]),
        .I2(\r7/t1/t0/p_0_in [3]),
        .I3(k6b[83]),
        .I4(\r7/t3/t2/p_1_in [3]),
        .I5(\r7/t3/t2/p_0_in [3]),
        .O(\r7/p_0_out [83]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[83]_i_1__6 
       (.I0(\r8/t0/t3/p_0_in [3]),
        .I1(\r8/t2/t1/p_1_in [3]),
        .I2(\r8/t1/t0/p_0_in [3]),
        .I3(k7b[83]),
        .I4(\r8/t3/t2/p_1_in [3]),
        .I5(\r8/t3/t2/p_0_in [3]),
        .O(\r8/p_0_out [83]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[83]_i_1__7 
       (.I0(\r9/t0/t3/p_0_in [3]),
        .I1(\r9/t2/t1/p_1_in [3]),
        .I2(\r9/t1/t0/p_0_in [3]),
        .I3(k8b[83]),
        .I4(\r9/t3/t2/p_1_in [3]),
        .I5(\r9/t3/t2/p_0_in [3]),
        .O(\r9/p_0_out [83]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair355" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[83]_i_1__8 
       (.I0(\a10/k1a [19]),
        .I1(\a10/k4a [19]),
        .I2(\rf/p_2_in [19]),
        .O(\rf/p_4_out [83]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[84]_i_1 
       (.I0(\r1/t0/t3/p_0_in [4]),
        .I1(\r1/t2/t1/p_1_in [4]),
        .I2(\r1/t1/t0/p_0_in [4]),
        .I3(k0b[84]),
        .I4(\r1/t3/t2/p_1_in [4]),
        .I5(\r1/t3/t2/p_0_in [4]),
        .O(\r1/p_0_out [84]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[84]_i_1__0 
       (.I0(\r2/t0/t3/p_0_in [4]),
        .I1(\r2/t2/t1/p_1_in [4]),
        .I2(\r2/t1/t0/p_0_in [4]),
        .I3(k1b[84]),
        .I4(\r2/t3/t2/p_1_in [4]),
        .I5(\r2/t3/t2/p_0_in [4]),
        .O(\r2/p_0_out [84]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[84]_i_1__1 
       (.I0(\r3/t0/t3/p_0_in [4]),
        .I1(\r3/t2/t1/p_1_in [4]),
        .I2(\r3/t1/t0/p_0_in [4]),
        .I3(k2b[84]),
        .I4(\r3/t3/t2/p_1_in [4]),
        .I5(\r3/t3/t2/p_0_in [4]),
        .O(\r3/p_0_out [84]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[84]_i_1__2 
       (.I0(\r4/t0/t3/p_0_in [4]),
        .I1(\r4/t2/t1/p_1_in [4]),
        .I2(\r4/t1/t0/p_0_in [4]),
        .I3(k3b[84]),
        .I4(\r4/t3/t2/p_1_in [4]),
        .I5(\r4/t3/t2/p_0_in [4]),
        .O(\r4/p_0_out [84]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[84]_i_1__3 
       (.I0(\r5/t0/t3/p_0_in [4]),
        .I1(\r5/t2/t1/p_1_in [4]),
        .I2(\r5/t1/t0/p_0_in [4]),
        .I3(k4b[84]),
        .I4(\r5/t3/t2/p_1_in [4]),
        .I5(\r5/t3/t2/p_0_in [4]),
        .O(\r5/p_0_out [84]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[84]_i_1__4 
       (.I0(\r6/t0/t3/p_0_in [4]),
        .I1(\r6/t2/t1/p_1_in [4]),
        .I2(\r6/t1/t0/p_0_in [4]),
        .I3(k5b[84]),
        .I4(\r6/t3/t2/p_1_in [4]),
        .I5(\r6/t3/t2/p_0_in [4]),
        .O(\r6/p_0_out [84]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[84]_i_1__5 
       (.I0(\r7/t0/t3/p_0_in [4]),
        .I1(\r7/t2/t1/p_1_in [4]),
        .I2(\r7/t1/t0/p_0_in [4]),
        .I3(k6b[84]),
        .I4(\r7/t3/t2/p_1_in [4]),
        .I5(\r7/t3/t2/p_0_in [4]),
        .O(\r7/p_0_out [84]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[84]_i_1__6 
       (.I0(\r8/t0/t3/p_0_in [4]),
        .I1(\r8/t2/t1/p_1_in [4]),
        .I2(\r8/t1/t0/p_0_in [4]),
        .I3(k7b[84]),
        .I4(\r8/t3/t2/p_1_in [4]),
        .I5(\r8/t3/t2/p_0_in [4]),
        .O(\r8/p_0_out [84]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[84]_i_1__7 
       (.I0(\r9/t0/t3/p_0_in [4]),
        .I1(\r9/t2/t1/p_1_in [4]),
        .I2(\r9/t1/t0/p_0_in [4]),
        .I3(k8b[84]),
        .I4(\r9/t3/t2/p_1_in [4]),
        .I5(\r9/t3/t2/p_0_in [4]),
        .O(\r9/p_0_out [84]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair354" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[84]_i_1__8 
       (.I0(\a10/k1a [20]),
        .I1(\a10/k4a [20]),
        .I2(\rf/p_2_in [20]),
        .O(\rf/p_4_out [84]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[85]_i_1 
       (.I0(\r1/t0/t3/p_0_in [5]),
        .I1(\r1/t2/t1/p_1_in [5]),
        .I2(\r1/t1/t0/p_0_in [5]),
        .I3(k0b[85]),
        .I4(\r1/t3/t2/p_1_in [5]),
        .I5(\r1/t3/t2/p_0_in [5]),
        .O(\r1/p_0_out [85]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[85]_i_1__0 
       (.I0(\r2/t0/t3/p_0_in [5]),
        .I1(\r2/t2/t1/p_1_in [5]),
        .I2(\r2/t1/t0/p_0_in [5]),
        .I3(k1b[85]),
        .I4(\r2/t3/t2/p_1_in [5]),
        .I5(\r2/t3/t2/p_0_in [5]),
        .O(\r2/p_0_out [85]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[85]_i_1__1 
       (.I0(\r3/t0/t3/p_0_in [5]),
        .I1(\r3/t2/t1/p_1_in [5]),
        .I2(\r3/t1/t0/p_0_in [5]),
        .I3(k2b[85]),
        .I4(\r3/t3/t2/p_1_in [5]),
        .I5(\r3/t3/t2/p_0_in [5]),
        .O(\r3/p_0_out [85]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[85]_i_1__2 
       (.I0(\r4/t0/t3/p_0_in [5]),
        .I1(\r4/t2/t1/p_1_in [5]),
        .I2(\r4/t1/t0/p_0_in [5]),
        .I3(k3b[85]),
        .I4(\r4/t3/t2/p_1_in [5]),
        .I5(\r4/t3/t2/p_0_in [5]),
        .O(\r4/p_0_out [85]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[85]_i_1__3 
       (.I0(\r5/t0/t3/p_0_in [5]),
        .I1(\r5/t2/t1/p_1_in [5]),
        .I2(\r5/t1/t0/p_0_in [5]),
        .I3(k4b[85]),
        .I4(\r5/t3/t2/p_1_in [5]),
        .I5(\r5/t3/t2/p_0_in [5]),
        .O(\r5/p_0_out [85]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[85]_i_1__4 
       (.I0(\r6/t0/t3/p_0_in [5]),
        .I1(\r6/t2/t1/p_1_in [5]),
        .I2(\r6/t1/t0/p_0_in [5]),
        .I3(k5b[85]),
        .I4(\r6/t3/t2/p_1_in [5]),
        .I5(\r6/t3/t2/p_0_in [5]),
        .O(\r6/p_0_out [85]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[85]_i_1__5 
       (.I0(\r7/t0/t3/p_0_in [5]),
        .I1(\r7/t2/t1/p_1_in [5]),
        .I2(\r7/t1/t0/p_0_in [5]),
        .I3(k6b[85]),
        .I4(\r7/t3/t2/p_1_in [5]),
        .I5(\r7/t3/t2/p_0_in [5]),
        .O(\r7/p_0_out [85]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[85]_i_1__6 
       (.I0(\r8/t0/t3/p_0_in [5]),
        .I1(\r8/t2/t1/p_1_in [5]),
        .I2(\r8/t1/t0/p_0_in [5]),
        .I3(k7b[85]),
        .I4(\r8/t3/t2/p_1_in [5]),
        .I5(\r8/t3/t2/p_0_in [5]),
        .O(\r8/p_0_out [85]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[85]_i_1__7 
       (.I0(\r9/t0/t3/p_0_in [5]),
        .I1(\r9/t2/t1/p_1_in [5]),
        .I2(\r9/t1/t0/p_0_in [5]),
        .I3(k8b[85]),
        .I4(\r9/t3/t2/p_1_in [5]),
        .I5(\r9/t3/t2/p_0_in [5]),
        .O(\r9/p_0_out [85]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair353" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[85]_i_1__8 
       (.I0(\a10/k1a [21]),
        .I1(\a10/k4a [21]),
        .I2(\rf/p_2_in [21]),
        .O(\rf/p_4_out [85]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[86]_i_1 
       (.I0(\r1/t0/t3/p_0_in [6]),
        .I1(\r1/t2/t1/p_1_in [6]),
        .I2(\r1/t1/t0/p_0_in [6]),
        .I3(k0b[86]),
        .I4(\r1/t3/t2/p_1_in [6]),
        .I5(\r1/t3/t2/p_0_in [6]),
        .O(\r1/p_0_out [86]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[86]_i_1__0 
       (.I0(\r2/t0/t3/p_0_in [6]),
        .I1(\r2/t2/t1/p_1_in [6]),
        .I2(\r2/t1/t0/p_0_in [6]),
        .I3(k1b[86]),
        .I4(\r2/t3/t2/p_1_in [6]),
        .I5(\r2/t3/t2/p_0_in [6]),
        .O(\r2/p_0_out [86]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[86]_i_1__1 
       (.I0(\r3/t0/t3/p_0_in [6]),
        .I1(\r3/t2/t1/p_1_in [6]),
        .I2(\r3/t1/t0/p_0_in [6]),
        .I3(k2b[86]),
        .I4(\r3/t3/t2/p_1_in [6]),
        .I5(\r3/t3/t2/p_0_in [6]),
        .O(\r3/p_0_out [86]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[86]_i_1__2 
       (.I0(\r4/t0/t3/p_0_in [6]),
        .I1(\r4/t2/t1/p_1_in [6]),
        .I2(\r4/t1/t0/p_0_in [6]),
        .I3(k3b[86]),
        .I4(\r4/t3/t2/p_1_in [6]),
        .I5(\r4/t3/t2/p_0_in [6]),
        .O(\r4/p_0_out [86]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[86]_i_1__3 
       (.I0(\r5/t0/t3/p_0_in [6]),
        .I1(\r5/t2/t1/p_1_in [6]),
        .I2(\r5/t1/t0/p_0_in [6]),
        .I3(k4b[86]),
        .I4(\r5/t3/t2/p_1_in [6]),
        .I5(\r5/t3/t2/p_0_in [6]),
        .O(\r5/p_0_out [86]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[86]_i_1__4 
       (.I0(\r6/t0/t3/p_0_in [6]),
        .I1(\r6/t2/t1/p_1_in [6]),
        .I2(\r6/t1/t0/p_0_in [6]),
        .I3(k5b[86]),
        .I4(\r6/t3/t2/p_1_in [6]),
        .I5(\r6/t3/t2/p_0_in [6]),
        .O(\r6/p_0_out [86]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[86]_i_1__5 
       (.I0(\r7/t0/t3/p_0_in [6]),
        .I1(\r7/t2/t1/p_1_in [6]),
        .I2(\r7/t1/t0/p_0_in [6]),
        .I3(k6b[86]),
        .I4(\r7/t3/t2/p_1_in [6]),
        .I5(\r7/t3/t2/p_0_in [6]),
        .O(\r7/p_0_out [86]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[86]_i_1__6 
       (.I0(\r8/t0/t3/p_0_in [6]),
        .I1(\r8/t2/t1/p_1_in [6]),
        .I2(\r8/t1/t0/p_0_in [6]),
        .I3(k7b[86]),
        .I4(\r8/t3/t2/p_1_in [6]),
        .I5(\r8/t3/t2/p_0_in [6]),
        .O(\r8/p_0_out [86]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[86]_i_1__7 
       (.I0(\r9/t0/t3/p_0_in [6]),
        .I1(\r9/t2/t1/p_1_in [6]),
        .I2(\r9/t1/t0/p_0_in [6]),
        .I3(k8b[86]),
        .I4(\r9/t3/t2/p_1_in [6]),
        .I5(\r9/t3/t2/p_0_in [6]),
        .O(\r9/p_0_out [86]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair352" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[86]_i_1__8 
       (.I0(\a10/k1a [22]),
        .I1(\a10/k4a [22]),
        .I2(\rf/p_2_in [22]),
        .O(\rf/p_4_out [86]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[87]_i_1 
       (.I0(\r1/t0/t3/p_0_in [7]),
        .I1(\r1/t2/t1/p_1_in [7]),
        .I2(\r1/t1/t0/p_0_in [7]),
        .I3(k0b[87]),
        .I4(\r1/t3/t2/p_1_in [7]),
        .I5(\r1/t3/t2/p_0_in [7]),
        .O(\r1/p_0_out [87]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[87]_i_1__0 
       (.I0(\r2/t0/t3/p_0_in [7]),
        .I1(\r2/t2/t1/p_1_in [7]),
        .I2(\r2/t1/t0/p_0_in [7]),
        .I3(k1b[87]),
        .I4(\r2/t3/t2/p_1_in [7]),
        .I5(\r2/t3/t2/p_0_in [7]),
        .O(\r2/p_0_out [87]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[87]_i_1__1 
       (.I0(\r3/t0/t3/p_0_in [7]),
        .I1(\r3/t2/t1/p_1_in [7]),
        .I2(\r3/t1/t0/p_0_in [7]),
        .I3(k2b[87]),
        .I4(\r3/t3/t2/p_1_in [7]),
        .I5(\r3/t3/t2/p_0_in [7]),
        .O(\r3/p_0_out [87]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[87]_i_1__2 
       (.I0(\r4/t0/t3/p_0_in [7]),
        .I1(\r4/t2/t1/p_1_in [7]),
        .I2(\r4/t1/t0/p_0_in [7]),
        .I3(k3b[87]),
        .I4(\r4/t3/t2/p_1_in [7]),
        .I5(\r4/t3/t2/p_0_in [7]),
        .O(\r4/p_0_out [87]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[87]_i_1__3 
       (.I0(\r5/t0/t3/p_0_in [7]),
        .I1(\r5/t2/t1/p_1_in [7]),
        .I2(\r5/t1/t0/p_0_in [7]),
        .I3(k4b[87]),
        .I4(\r5/t3/t2/p_1_in [7]),
        .I5(\r5/t3/t2/p_0_in [7]),
        .O(\r5/p_0_out [87]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[87]_i_1__4 
       (.I0(\r6/t0/t3/p_0_in [7]),
        .I1(\r6/t2/t1/p_1_in [7]),
        .I2(\r6/t1/t0/p_0_in [7]),
        .I3(k5b[87]),
        .I4(\r6/t3/t2/p_1_in [7]),
        .I5(\r6/t3/t2/p_0_in [7]),
        .O(\r6/p_0_out [87]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[87]_i_1__5 
       (.I0(\r7/t0/t3/p_0_in [7]),
        .I1(\r7/t2/t1/p_1_in [7]),
        .I2(\r7/t1/t0/p_0_in [7]),
        .I3(k6b[87]),
        .I4(\r7/t3/t2/p_1_in [7]),
        .I5(\r7/t3/t2/p_0_in [7]),
        .O(\r7/p_0_out [87]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[87]_i_1__6 
       (.I0(\r8/t0/t3/p_0_in [7]),
        .I1(\r8/t2/t1/p_1_in [7]),
        .I2(\r8/t1/t0/p_0_in [7]),
        .I3(k7b[87]),
        .I4(\r8/t3/t2/p_1_in [7]),
        .I5(\r8/t3/t2/p_0_in [7]),
        .O(\r8/p_0_out [87]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[87]_i_1__7 
       (.I0(\r9/t0/t3/p_0_in [7]),
        .I1(\r9/t2/t1/p_1_in [7]),
        .I2(\r9/t1/t0/p_0_in [7]),
        .I3(k8b[87]),
        .I4(\r9/t3/t2/p_1_in [7]),
        .I5(\r9/t3/t2/p_0_in [7]),
        .O(\r9/p_0_out [87]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair351" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[87]_i_1__8 
       (.I0(\a10/k1a [23]),
        .I1(\a10/k4a [23]),
        .I2(\rf/p_2_in [23]),
        .O(\rf/p_4_out [87]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[88]_i_1 
       (.I0(\r1/t0/t3/p_0_in [0]),
        .I1(\r1/t2/t1/p_1_in [0]),
        .I2(\r1/t2/t1/p_0_in [0]),
        .I3(\r1/t1/t0/p_1_in [0]),
        .I4(k0b[88]),
        .I5(\r1/t3/t2/p_0_in [0]),
        .O(\r1/p_0_out [88]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[88]_i_1__0 
       (.I0(\r2/t0/t3/p_0_in [0]),
        .I1(\r2/t2/t1/p_1_in [0]),
        .I2(\r2/t2/t1/p_0_in [0]),
        .I3(\r2/t1/t0/p_1_in [0]),
        .I4(k1b[88]),
        .I5(\r2/t3/t2/p_0_in [0]),
        .O(\r2/p_0_out [88]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[88]_i_1__1 
       (.I0(\r3/t0/t3/p_0_in [0]),
        .I1(\r3/t2/t1/p_1_in [0]),
        .I2(\r3/t2/t1/p_0_in [0]),
        .I3(\r3/t1/t0/p_1_in [0]),
        .I4(k2b[88]),
        .I5(\r3/t3/t2/p_0_in [0]),
        .O(\r3/p_0_out [88]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[88]_i_1__2 
       (.I0(\r4/t0/t3/p_0_in [0]),
        .I1(\r4/t2/t1/p_1_in [0]),
        .I2(\r4/t2/t1/p_0_in [0]),
        .I3(\r4/t1/t0/p_1_in [0]),
        .I4(k3b[88]),
        .I5(\r4/t3/t2/p_0_in [0]),
        .O(\r4/p_0_out [88]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[88]_i_1__3 
       (.I0(\r5/t0/t3/p_0_in [0]),
        .I1(\r5/t2/t1/p_1_in [0]),
        .I2(\r5/t2/t1/p_0_in [0]),
        .I3(\r5/t1/t0/p_1_in [0]),
        .I4(k4b[88]),
        .I5(\r5/t3/t2/p_0_in [0]),
        .O(\r5/p_0_out [88]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[88]_i_1__4 
       (.I0(\r6/t0/t3/p_0_in [0]),
        .I1(\r6/t2/t1/p_1_in [0]),
        .I2(\r6/t2/t1/p_0_in [0]),
        .I3(\r6/t1/t0/p_1_in [0]),
        .I4(k5b[88]),
        .I5(\r6/t3/t2/p_0_in [0]),
        .O(\r6/p_0_out [88]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[88]_i_1__5 
       (.I0(\r7/t0/t3/p_0_in [0]),
        .I1(\r7/t2/t1/p_1_in [0]),
        .I2(\r7/t2/t1/p_0_in [0]),
        .I3(\r7/t1/t0/p_1_in [0]),
        .I4(k6b[88]),
        .I5(\r7/t3/t2/p_0_in [0]),
        .O(\r7/p_0_out [88]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[88]_i_1__6 
       (.I0(\r8/t0/t3/p_0_in [0]),
        .I1(\r8/t2/t1/p_1_in [0]),
        .I2(\r8/t2/t1/p_0_in [0]),
        .I3(\r8/t1/t0/p_1_in [0]),
        .I4(k7b[88]),
        .I5(\r8/t3/t2/p_0_in [0]),
        .O(\r8/p_0_out [88]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[88]_i_1__7 
       (.I0(\r9/t0/t3/p_0_in [0]),
        .I1(\r9/t2/t1/p_1_in [0]),
        .I2(\r9/t2/t1/p_0_in [0]),
        .I3(\r9/t1/t0/p_1_in [0]),
        .I4(k8b[88]),
        .I5(\r9/t3/t2/p_0_in [0]),
        .O(\r9/p_0_out [88]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair350" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[88]_i_1__8 
       (.I0(\a10/k1a [24]),
        .I1(\a10/k4a [24]),
        .I2(\rf/p_2_in [24]),
        .O(\rf/p_4_out [88]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[89]_i_1 
       (.I0(\r1/t0/t3/p_0_in [1]),
        .I1(\r1/t2/t1/p_1_in [1]),
        .I2(\r1/t2/t1/p_0_in [1]),
        .I3(\r1/t1/t0/p_1_in [1]),
        .I4(k0b[89]),
        .I5(\r1/t3/t2/p_0_in [1]),
        .O(\r1/p_0_out [89]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[89]_i_1__0 
       (.I0(\r2/t0/t3/p_0_in [1]),
        .I1(\r2/t2/t1/p_1_in [1]),
        .I2(\r2/t2/t1/p_0_in [1]),
        .I3(\r2/t1/t0/p_1_in [1]),
        .I4(k1b[89]),
        .I5(\r2/t3/t2/p_0_in [1]),
        .O(\r2/p_0_out [89]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[89]_i_1__1 
       (.I0(\r3/t0/t3/p_0_in [1]),
        .I1(\r3/t2/t1/p_1_in [1]),
        .I2(\r3/t2/t1/p_0_in [1]),
        .I3(\r3/t1/t0/p_1_in [1]),
        .I4(k2b[89]),
        .I5(\r3/t3/t2/p_0_in [1]),
        .O(\r3/p_0_out [89]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[89]_i_1__2 
       (.I0(\r4/t0/t3/p_0_in [1]),
        .I1(\r4/t2/t1/p_1_in [1]),
        .I2(\r4/t2/t1/p_0_in [1]),
        .I3(\r4/t1/t0/p_1_in [1]),
        .I4(k3b[89]),
        .I5(\r4/t3/t2/p_0_in [1]),
        .O(\r4/p_0_out [89]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[89]_i_1__3 
       (.I0(\r5/t0/t3/p_0_in [1]),
        .I1(\r5/t2/t1/p_1_in [1]),
        .I2(\r5/t2/t1/p_0_in [1]),
        .I3(\r5/t1/t0/p_1_in [1]),
        .I4(k4b[89]),
        .I5(\r5/t3/t2/p_0_in [1]),
        .O(\r5/p_0_out [89]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[89]_i_1__4 
       (.I0(\r6/t0/t3/p_0_in [1]),
        .I1(\r6/t2/t1/p_1_in [1]),
        .I2(\r6/t2/t1/p_0_in [1]),
        .I3(\r6/t1/t0/p_1_in [1]),
        .I4(k5b[89]),
        .I5(\r6/t3/t2/p_0_in [1]),
        .O(\r6/p_0_out [89]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[89]_i_1__5 
       (.I0(\r7/t0/t3/p_0_in [1]),
        .I1(\r7/t2/t1/p_1_in [1]),
        .I2(\r7/t2/t1/p_0_in [1]),
        .I3(\r7/t1/t0/p_1_in [1]),
        .I4(k6b[89]),
        .I5(\r7/t3/t2/p_0_in [1]),
        .O(\r7/p_0_out [89]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[89]_i_1__6 
       (.I0(\r8/t0/t3/p_0_in [1]),
        .I1(\r8/t2/t1/p_1_in [1]),
        .I2(\r8/t2/t1/p_0_in [1]),
        .I3(\r8/t1/t0/p_1_in [1]),
        .I4(k7b[89]),
        .I5(\r8/t3/t2/p_0_in [1]),
        .O(\r8/p_0_out [89]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[89]_i_1__7 
       (.I0(\r9/t0/t3/p_0_in [1]),
        .I1(\r9/t2/t1/p_1_in [1]),
        .I2(\r9/t2/t1/p_0_in [1]),
        .I3(\r9/t1/t0/p_1_in [1]),
        .I4(k8b[89]),
        .I5(\r9/t3/t2/p_0_in [1]),
        .O(\r9/p_0_out [89]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair349" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[89]_i_1__8 
       (.I0(\a10/k1a [25]),
        .I1(\a10/k4a [25]),
        .I2(\rf/p_2_in [25]),
        .O(\rf/p_4_out [89]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[8]_i_1 
       (.I0(\r1/t0/t1/p_0_in [0]),
        .I1(\r1/t2/t3/p_1_in [0]),
        .I2(\r1/t2/t3/p_0_in [0]),
        .I3(\r1/t1/t2/p_1_in [0]),
        .I4(k0b[8]),
        .I5(\r1/t3/t0/p_0_in [0]),
        .O(\r1/p_0_out [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[8]_i_1__0 
       (.I0(\r2/t0/t1/p_0_in [0]),
        .I1(\r2/t2/t3/p_1_in [0]),
        .I2(\r2/t2/t3/p_0_in [0]),
        .I3(\r2/t1/t2/p_1_in [0]),
        .I4(k1b[8]),
        .I5(\r2/t3/t0/p_0_in [0]),
        .O(\r2/p_0_out [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[8]_i_1__1 
       (.I0(\r3/t0/t1/p_0_in [0]),
        .I1(\r3/t2/t3/p_1_in [0]),
        .I2(\r3/t2/t3/p_0_in [0]),
        .I3(\r3/t1/t2/p_1_in [0]),
        .I4(k2b[8]),
        .I5(\r3/t3/t0/p_0_in [0]),
        .O(\r3/p_0_out [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[8]_i_1__2 
       (.I0(\r4/t0/t1/p_0_in [0]),
        .I1(\r4/t2/t3/p_1_in [0]),
        .I2(\r4/t2/t3/p_0_in [0]),
        .I3(\r4/t1/t2/p_1_in [0]),
        .I4(k3b[8]),
        .I5(\r4/t3/t0/p_0_in [0]),
        .O(\r4/p_0_out [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[8]_i_1__3 
       (.I0(\r5/t0/t1/p_0_in [0]),
        .I1(\r5/t2/t3/p_1_in [0]),
        .I2(\r5/t2/t3/p_0_in [0]),
        .I3(\r5/t1/t2/p_1_in [0]),
        .I4(k4b[8]),
        .I5(\r5/t3/t0/p_0_in [0]),
        .O(\r5/p_0_out [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[8]_i_1__4 
       (.I0(\r6/t0/t1/p_0_in [0]),
        .I1(\r6/t2/t3/p_1_in [0]),
        .I2(\r6/t2/t3/p_0_in [0]),
        .I3(\r6/t1/t2/p_1_in [0]),
        .I4(k5b[8]),
        .I5(\r6/t3/t0/p_0_in [0]),
        .O(\r6/p_0_out [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[8]_i_1__5 
       (.I0(\r7/t0/t1/p_0_in [0]),
        .I1(\r7/t2/t3/p_1_in [0]),
        .I2(\r7/t2/t3/p_0_in [0]),
        .I3(\r7/t1/t2/p_1_in [0]),
        .I4(k6b[8]),
        .I5(\r7/t3/t0/p_0_in [0]),
        .O(\r7/p_0_out [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[8]_i_1__6 
       (.I0(\r8/t0/t1/p_0_in [0]),
        .I1(\r8/t2/t3/p_1_in [0]),
        .I2(\r8/t2/t3/p_0_in [0]),
        .I3(\r8/t1/t2/p_1_in [0]),
        .I4(k7b[8]),
        .I5(\r8/t3/t0/p_0_in [0]),
        .O(\r8/p_0_out [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[8]_i_1__7 
       (.I0(\r9/t0/t1/p_0_in [0]),
        .I1(\r9/t2/t3/p_1_in [0]),
        .I2(\r9/t2/t3/p_0_in [0]),
        .I3(\r9/t1/t2/p_1_in [0]),
        .I4(k8b[8]),
        .I5(\r9/t3/t0/p_0_in [0]),
        .O(\r9/p_0_out [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair334" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[8]_i_1__8 
       (.I0(\a10/k3a [8]),
        .I1(\a10/k4a [8]),
        .I2(\rf/p_0_in [8]),
        .O(\rf/p_4_out [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[90]_i_1 
       (.I0(\r1/t0/t3/p_0_in [2]),
        .I1(\r1/t2/t1/p_1_in [2]),
        .I2(\r1/t2/t1/p_0_in [2]),
        .I3(\r1/t1/t0/p_1_in [2]),
        .I4(k0b[90]),
        .I5(\r1/t3/t2/p_0_in [2]),
        .O(\r1/p_0_out [90]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[90]_i_1__0 
       (.I0(\r2/t0/t3/p_0_in [2]),
        .I1(\r2/t2/t1/p_1_in [2]),
        .I2(\r2/t2/t1/p_0_in [2]),
        .I3(\r2/t1/t0/p_1_in [2]),
        .I4(k1b[90]),
        .I5(\r2/t3/t2/p_0_in [2]),
        .O(\r2/p_0_out [90]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[90]_i_1__1 
       (.I0(\r3/t0/t3/p_0_in [2]),
        .I1(\r3/t2/t1/p_1_in [2]),
        .I2(\r3/t2/t1/p_0_in [2]),
        .I3(\r3/t1/t0/p_1_in [2]),
        .I4(k2b[90]),
        .I5(\r3/t3/t2/p_0_in [2]),
        .O(\r3/p_0_out [90]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[90]_i_1__2 
       (.I0(\r4/t0/t3/p_0_in [2]),
        .I1(\r4/t2/t1/p_1_in [2]),
        .I2(\r4/t2/t1/p_0_in [2]),
        .I3(\r4/t1/t0/p_1_in [2]),
        .I4(k3b[90]),
        .I5(\r4/t3/t2/p_0_in [2]),
        .O(\r4/p_0_out [90]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[90]_i_1__3 
       (.I0(\r5/t0/t3/p_0_in [2]),
        .I1(\r5/t2/t1/p_1_in [2]),
        .I2(\r5/t2/t1/p_0_in [2]),
        .I3(\r5/t1/t0/p_1_in [2]),
        .I4(k4b[90]),
        .I5(\r5/t3/t2/p_0_in [2]),
        .O(\r5/p_0_out [90]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[90]_i_1__4 
       (.I0(\r6/t0/t3/p_0_in [2]),
        .I1(\r6/t2/t1/p_1_in [2]),
        .I2(\r6/t2/t1/p_0_in [2]),
        .I3(\r6/t1/t0/p_1_in [2]),
        .I4(k5b[90]),
        .I5(\r6/t3/t2/p_0_in [2]),
        .O(\r6/p_0_out [90]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[90]_i_1__5 
       (.I0(\r7/t0/t3/p_0_in [2]),
        .I1(\r7/t2/t1/p_1_in [2]),
        .I2(\r7/t2/t1/p_0_in [2]),
        .I3(\r7/t1/t0/p_1_in [2]),
        .I4(k6b[90]),
        .I5(\r7/t3/t2/p_0_in [2]),
        .O(\r7/p_0_out [90]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[90]_i_1__6 
       (.I0(\r8/t0/t3/p_0_in [2]),
        .I1(\r8/t2/t1/p_1_in [2]),
        .I2(\r8/t2/t1/p_0_in [2]),
        .I3(\r8/t1/t0/p_1_in [2]),
        .I4(k7b[90]),
        .I5(\r8/t3/t2/p_0_in [2]),
        .O(\r8/p_0_out [90]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[90]_i_1__7 
       (.I0(\r9/t0/t3/p_0_in [2]),
        .I1(\r9/t2/t1/p_1_in [2]),
        .I2(\r9/t2/t1/p_0_in [2]),
        .I3(\r9/t1/t0/p_1_in [2]),
        .I4(k8b[90]),
        .I5(\r9/t3/t2/p_0_in [2]),
        .O(\r9/p_0_out [90]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair348" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[90]_i_1__8 
       (.I0(\a10/k1a [26]),
        .I1(\a10/k4a [26]),
        .I2(\rf/p_2_in [26]),
        .O(\rf/p_4_out [90]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[91]_i_1 
       (.I0(\r1/t0/t3/p_0_in [3]),
        .I1(\r1/t2/t1/p_1_in [3]),
        .I2(\r1/t2/t1/p_0_in [3]),
        .I3(\r1/t1/t0/p_1_in [3]),
        .I4(k0b[91]),
        .I5(\r1/t3/t2/p_0_in [3]),
        .O(\r1/p_0_out [91]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[91]_i_1__0 
       (.I0(\r2/t0/t3/p_0_in [3]),
        .I1(\r2/t2/t1/p_1_in [3]),
        .I2(\r2/t2/t1/p_0_in [3]),
        .I3(\r2/t1/t0/p_1_in [3]),
        .I4(k1b[91]),
        .I5(\r2/t3/t2/p_0_in [3]),
        .O(\r2/p_0_out [91]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[91]_i_1__1 
       (.I0(\r3/t0/t3/p_0_in [3]),
        .I1(\r3/t2/t1/p_1_in [3]),
        .I2(\r3/t2/t1/p_0_in [3]),
        .I3(\r3/t1/t0/p_1_in [3]),
        .I4(k2b[91]),
        .I5(\r3/t3/t2/p_0_in [3]),
        .O(\r3/p_0_out [91]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[91]_i_1__2 
       (.I0(\r4/t0/t3/p_0_in [3]),
        .I1(\r4/t2/t1/p_1_in [3]),
        .I2(\r4/t2/t1/p_0_in [3]),
        .I3(\r4/t1/t0/p_1_in [3]),
        .I4(k3b[91]),
        .I5(\r4/t3/t2/p_0_in [3]),
        .O(\r4/p_0_out [91]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[91]_i_1__3 
       (.I0(\r5/t0/t3/p_0_in [3]),
        .I1(\r5/t2/t1/p_1_in [3]),
        .I2(\r5/t2/t1/p_0_in [3]),
        .I3(\r5/t1/t0/p_1_in [3]),
        .I4(k4b[91]),
        .I5(\r5/t3/t2/p_0_in [3]),
        .O(\r5/p_0_out [91]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[91]_i_1__4 
       (.I0(\r6/t0/t3/p_0_in [3]),
        .I1(\r6/t2/t1/p_1_in [3]),
        .I2(\r6/t2/t1/p_0_in [3]),
        .I3(\r6/t1/t0/p_1_in [3]),
        .I4(k5b[91]),
        .I5(\r6/t3/t2/p_0_in [3]),
        .O(\r6/p_0_out [91]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[91]_i_1__5 
       (.I0(\r7/t0/t3/p_0_in [3]),
        .I1(\r7/t2/t1/p_1_in [3]),
        .I2(\r7/t2/t1/p_0_in [3]),
        .I3(\r7/t1/t0/p_1_in [3]),
        .I4(k6b[91]),
        .I5(\r7/t3/t2/p_0_in [3]),
        .O(\r7/p_0_out [91]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[91]_i_1__6 
       (.I0(\r8/t0/t3/p_0_in [3]),
        .I1(\r8/t2/t1/p_1_in [3]),
        .I2(\r8/t2/t1/p_0_in [3]),
        .I3(\r8/t1/t0/p_1_in [3]),
        .I4(k7b[91]),
        .I5(\r8/t3/t2/p_0_in [3]),
        .O(\r8/p_0_out [91]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[91]_i_1__7 
       (.I0(\r9/t0/t3/p_0_in [3]),
        .I1(\r9/t2/t1/p_1_in [3]),
        .I2(\r9/t2/t1/p_0_in [3]),
        .I3(\r9/t1/t0/p_1_in [3]),
        .I4(k8b[91]),
        .I5(\r9/t3/t2/p_0_in [3]),
        .O(\r9/p_0_out [91]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair347" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[91]_i_1__8 
       (.I0(\a10/k1a [27]),
        .I1(\a10/k4a [27]),
        .I2(\rf/p_2_in [27]),
        .O(\rf/p_4_out [91]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[92]_i_1 
       (.I0(\r1/t0/t3/p_0_in [4]),
        .I1(\r1/t2/t1/p_1_in [4]),
        .I2(\r1/t2/t1/p_0_in [4]),
        .I3(\r1/t1/t0/p_1_in [4]),
        .I4(k0b[92]),
        .I5(\r1/t3/t2/p_0_in [4]),
        .O(\r1/p_0_out [92]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[92]_i_1__0 
       (.I0(\r2/t0/t3/p_0_in [4]),
        .I1(\r2/t2/t1/p_1_in [4]),
        .I2(\r2/t2/t1/p_0_in [4]),
        .I3(\r2/t1/t0/p_1_in [4]),
        .I4(k1b[92]),
        .I5(\r2/t3/t2/p_0_in [4]),
        .O(\r2/p_0_out [92]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[92]_i_1__1 
       (.I0(\r3/t0/t3/p_0_in [4]),
        .I1(\r3/t2/t1/p_1_in [4]),
        .I2(\r3/t2/t1/p_0_in [4]),
        .I3(\r3/t1/t0/p_1_in [4]),
        .I4(k2b[92]),
        .I5(\r3/t3/t2/p_0_in [4]),
        .O(\r3/p_0_out [92]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[92]_i_1__2 
       (.I0(\r4/t0/t3/p_0_in [4]),
        .I1(\r4/t2/t1/p_1_in [4]),
        .I2(\r4/t2/t1/p_0_in [4]),
        .I3(\r4/t1/t0/p_1_in [4]),
        .I4(k3b[92]),
        .I5(\r4/t3/t2/p_0_in [4]),
        .O(\r4/p_0_out [92]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[92]_i_1__3 
       (.I0(\r5/t0/t3/p_0_in [4]),
        .I1(\r5/t2/t1/p_1_in [4]),
        .I2(\r5/t2/t1/p_0_in [4]),
        .I3(\r5/t1/t0/p_1_in [4]),
        .I4(k4b[92]),
        .I5(\r5/t3/t2/p_0_in [4]),
        .O(\r5/p_0_out [92]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[92]_i_1__4 
       (.I0(\r6/t0/t3/p_0_in [4]),
        .I1(\r6/t2/t1/p_1_in [4]),
        .I2(\r6/t2/t1/p_0_in [4]),
        .I3(\r6/t1/t0/p_1_in [4]),
        .I4(k5b[92]),
        .I5(\r6/t3/t2/p_0_in [4]),
        .O(\r6/p_0_out [92]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[92]_i_1__5 
       (.I0(\r7/t0/t3/p_0_in [4]),
        .I1(\r7/t2/t1/p_1_in [4]),
        .I2(\r7/t2/t1/p_0_in [4]),
        .I3(\r7/t1/t0/p_1_in [4]),
        .I4(k6b[92]),
        .I5(\r7/t3/t2/p_0_in [4]),
        .O(\r7/p_0_out [92]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[92]_i_1__6 
       (.I0(\r8/t0/t3/p_0_in [4]),
        .I1(\r8/t2/t1/p_1_in [4]),
        .I2(\r8/t2/t1/p_0_in [4]),
        .I3(\r8/t1/t0/p_1_in [4]),
        .I4(k7b[92]),
        .I5(\r8/t3/t2/p_0_in [4]),
        .O(\r8/p_0_out [92]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[92]_i_1__7 
       (.I0(\r9/t0/t3/p_0_in [4]),
        .I1(\r9/t2/t1/p_1_in [4]),
        .I2(\r9/t2/t1/p_0_in [4]),
        .I3(\r9/t1/t0/p_1_in [4]),
        .I4(k8b[92]),
        .I5(\r9/t3/t2/p_0_in [4]),
        .O(\r9/p_0_out [92]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair346" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[92]_i_1__8 
       (.I0(\a10/k1a [28]),
        .I1(\a10/k4a [28]),
        .I2(\rf/p_2_in [28]),
        .O(\rf/p_4_out [92]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[93]_i_1 
       (.I0(\r1/t0/t3/p_0_in [5]),
        .I1(\r1/t2/t1/p_1_in [5]),
        .I2(\r1/t2/t1/p_0_in [5]),
        .I3(\r1/t1/t0/p_1_in [5]),
        .I4(k0b[93]),
        .I5(\r1/t3/t2/p_0_in [5]),
        .O(\r1/p_0_out [93]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[93]_i_1__0 
       (.I0(\r2/t0/t3/p_0_in [5]),
        .I1(\r2/t2/t1/p_1_in [5]),
        .I2(\r2/t2/t1/p_0_in [5]),
        .I3(\r2/t1/t0/p_1_in [5]),
        .I4(k1b[93]),
        .I5(\r2/t3/t2/p_0_in [5]),
        .O(\r2/p_0_out [93]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[93]_i_1__1 
       (.I0(\r3/t0/t3/p_0_in [5]),
        .I1(\r3/t2/t1/p_1_in [5]),
        .I2(\r3/t2/t1/p_0_in [5]),
        .I3(\r3/t1/t0/p_1_in [5]),
        .I4(k2b[93]),
        .I5(\r3/t3/t2/p_0_in [5]),
        .O(\r3/p_0_out [93]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[93]_i_1__2 
       (.I0(\r4/t0/t3/p_0_in [5]),
        .I1(\r4/t2/t1/p_1_in [5]),
        .I2(\r4/t2/t1/p_0_in [5]),
        .I3(\r4/t1/t0/p_1_in [5]),
        .I4(k3b[93]),
        .I5(\r4/t3/t2/p_0_in [5]),
        .O(\r4/p_0_out [93]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[93]_i_1__3 
       (.I0(\r5/t0/t3/p_0_in [5]),
        .I1(\r5/t2/t1/p_1_in [5]),
        .I2(\r5/t2/t1/p_0_in [5]),
        .I3(\r5/t1/t0/p_1_in [5]),
        .I4(k4b[93]),
        .I5(\r5/t3/t2/p_0_in [5]),
        .O(\r5/p_0_out [93]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[93]_i_1__4 
       (.I0(\r6/t0/t3/p_0_in [5]),
        .I1(\r6/t2/t1/p_1_in [5]),
        .I2(\r6/t2/t1/p_0_in [5]),
        .I3(\r6/t1/t0/p_1_in [5]),
        .I4(k5b[93]),
        .I5(\r6/t3/t2/p_0_in [5]),
        .O(\r6/p_0_out [93]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[93]_i_1__5 
       (.I0(\r7/t0/t3/p_0_in [5]),
        .I1(\r7/t2/t1/p_1_in [5]),
        .I2(\r7/t2/t1/p_0_in [5]),
        .I3(\r7/t1/t0/p_1_in [5]),
        .I4(k6b[93]),
        .I5(\r7/t3/t2/p_0_in [5]),
        .O(\r7/p_0_out [93]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[93]_i_1__6 
       (.I0(\r8/t0/t3/p_0_in [5]),
        .I1(\r8/t2/t1/p_1_in [5]),
        .I2(\r8/t2/t1/p_0_in [5]),
        .I3(\r8/t1/t0/p_1_in [5]),
        .I4(k7b[93]),
        .I5(\r8/t3/t2/p_0_in [5]),
        .O(\r8/p_0_out [93]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[93]_i_1__7 
       (.I0(\r9/t0/t3/p_0_in [5]),
        .I1(\r9/t2/t1/p_1_in [5]),
        .I2(\r9/t2/t1/p_0_in [5]),
        .I3(\r9/t1/t0/p_1_in [5]),
        .I4(k8b[93]),
        .I5(\r9/t3/t2/p_0_in [5]),
        .O(\r9/p_0_out [93]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair345" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[93]_i_1__8 
       (.I0(\a10/k1a [29]),
        .I1(\a10/k4a [29]),
        .I2(\rf/p_2_in [29]),
        .O(\rf/p_4_out [93]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[94]_i_1 
       (.I0(\r1/t0/t3/p_0_in [6]),
        .I1(\r1/t2/t1/p_1_in [6]),
        .I2(\r1/t2/t1/p_0_in [6]),
        .I3(\r1/t1/t0/p_1_in [6]),
        .I4(k0b[94]),
        .I5(\r1/t3/t2/p_0_in [6]),
        .O(\r1/p_0_out [94]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[94]_i_1__0 
       (.I0(\r2/t0/t3/p_0_in [6]),
        .I1(\r2/t2/t1/p_1_in [6]),
        .I2(\r2/t2/t1/p_0_in [6]),
        .I3(\r2/t1/t0/p_1_in [6]),
        .I4(k1b[94]),
        .I5(\r2/t3/t2/p_0_in [6]),
        .O(\r2/p_0_out [94]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[94]_i_1__1 
       (.I0(\r3/t0/t3/p_0_in [6]),
        .I1(\r3/t2/t1/p_1_in [6]),
        .I2(\r3/t2/t1/p_0_in [6]),
        .I3(\r3/t1/t0/p_1_in [6]),
        .I4(k2b[94]),
        .I5(\r3/t3/t2/p_0_in [6]),
        .O(\r3/p_0_out [94]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[94]_i_1__2 
       (.I0(\r4/t0/t3/p_0_in [6]),
        .I1(\r4/t2/t1/p_1_in [6]),
        .I2(\r4/t2/t1/p_0_in [6]),
        .I3(\r4/t1/t0/p_1_in [6]),
        .I4(k3b[94]),
        .I5(\r4/t3/t2/p_0_in [6]),
        .O(\r4/p_0_out [94]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[94]_i_1__3 
       (.I0(\r5/t0/t3/p_0_in [6]),
        .I1(\r5/t2/t1/p_1_in [6]),
        .I2(\r5/t2/t1/p_0_in [6]),
        .I3(\r5/t1/t0/p_1_in [6]),
        .I4(k4b[94]),
        .I5(\r5/t3/t2/p_0_in [6]),
        .O(\r5/p_0_out [94]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[94]_i_1__4 
       (.I0(\r6/t0/t3/p_0_in [6]),
        .I1(\r6/t2/t1/p_1_in [6]),
        .I2(\r6/t2/t1/p_0_in [6]),
        .I3(\r6/t1/t0/p_1_in [6]),
        .I4(k5b[94]),
        .I5(\r6/t3/t2/p_0_in [6]),
        .O(\r6/p_0_out [94]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[94]_i_1__5 
       (.I0(\r7/t0/t3/p_0_in [6]),
        .I1(\r7/t2/t1/p_1_in [6]),
        .I2(\r7/t2/t1/p_0_in [6]),
        .I3(\r7/t1/t0/p_1_in [6]),
        .I4(k6b[94]),
        .I5(\r7/t3/t2/p_0_in [6]),
        .O(\r7/p_0_out [94]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[94]_i_1__6 
       (.I0(\r8/t0/t3/p_0_in [6]),
        .I1(\r8/t2/t1/p_1_in [6]),
        .I2(\r8/t2/t1/p_0_in [6]),
        .I3(\r8/t1/t0/p_1_in [6]),
        .I4(k7b[94]),
        .I5(\r8/t3/t2/p_0_in [6]),
        .O(\r8/p_0_out [94]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[94]_i_1__7 
       (.I0(\r9/t0/t3/p_0_in [6]),
        .I1(\r9/t2/t1/p_1_in [6]),
        .I2(\r9/t2/t1/p_0_in [6]),
        .I3(\r9/t1/t0/p_1_in [6]),
        .I4(k8b[94]),
        .I5(\r9/t3/t2/p_0_in [6]),
        .O(\r9/p_0_out [94]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair344" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[94]_i_1__8 
       (.I0(\a10/k1a [30]),
        .I1(\a10/k4a [30]),
        .I2(\rf/p_2_in [30]),
        .O(\rf/p_4_out [94]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[95]_i_1 
       (.I0(\r1/t0/t3/p_0_in [7]),
        .I1(\r1/t2/t1/p_1_in [7]),
        .I2(\r1/t2/t1/p_0_in [7]),
        .I3(\r1/t1/t0/p_1_in [7]),
        .I4(k0b[95]),
        .I5(\r1/t3/t2/p_0_in [7]),
        .O(\r1/p_0_out [95]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[95]_i_1__0 
       (.I0(\r2/t0/t3/p_0_in [7]),
        .I1(\r2/t2/t1/p_1_in [7]),
        .I2(\r2/t2/t1/p_0_in [7]),
        .I3(\r2/t1/t0/p_1_in [7]),
        .I4(k1b[95]),
        .I5(\r2/t3/t2/p_0_in [7]),
        .O(\r2/p_0_out [95]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[95]_i_1__1 
       (.I0(\r3/t0/t3/p_0_in [7]),
        .I1(\r3/t2/t1/p_1_in [7]),
        .I2(\r3/t2/t1/p_0_in [7]),
        .I3(\r3/t1/t0/p_1_in [7]),
        .I4(k2b[95]),
        .I5(\r3/t3/t2/p_0_in [7]),
        .O(\r3/p_0_out [95]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[95]_i_1__2 
       (.I0(\r4/t0/t3/p_0_in [7]),
        .I1(\r4/t2/t1/p_1_in [7]),
        .I2(\r4/t2/t1/p_0_in [7]),
        .I3(\r4/t1/t0/p_1_in [7]),
        .I4(k3b[95]),
        .I5(\r4/t3/t2/p_0_in [7]),
        .O(\r4/p_0_out [95]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[95]_i_1__3 
       (.I0(\r5/t0/t3/p_0_in [7]),
        .I1(\r5/t2/t1/p_1_in [7]),
        .I2(\r5/t2/t1/p_0_in [7]),
        .I3(\r5/t1/t0/p_1_in [7]),
        .I4(k4b[95]),
        .I5(\r5/t3/t2/p_0_in [7]),
        .O(\r5/p_0_out [95]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[95]_i_1__4 
       (.I0(\r6/t0/t3/p_0_in [7]),
        .I1(\r6/t2/t1/p_1_in [7]),
        .I2(\r6/t2/t1/p_0_in [7]),
        .I3(\r6/t1/t0/p_1_in [7]),
        .I4(k5b[95]),
        .I5(\r6/t3/t2/p_0_in [7]),
        .O(\r6/p_0_out [95]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[95]_i_1__5 
       (.I0(\r7/t0/t3/p_0_in [7]),
        .I1(\r7/t2/t1/p_1_in [7]),
        .I2(\r7/t2/t1/p_0_in [7]),
        .I3(\r7/t1/t0/p_1_in [7]),
        .I4(k6b[95]),
        .I5(\r7/t3/t2/p_0_in [7]),
        .O(\r7/p_0_out [95]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[95]_i_1__6 
       (.I0(\r8/t0/t3/p_0_in [7]),
        .I1(\r8/t2/t1/p_1_in [7]),
        .I2(\r8/t2/t1/p_0_in [7]),
        .I3(\r8/t1/t0/p_1_in [7]),
        .I4(k7b[95]),
        .I5(\r8/t3/t2/p_0_in [7]),
        .O(\r8/p_0_out [95]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[95]_i_1__7 
       (.I0(\r9/t0/t3/p_0_in [7]),
        .I1(\r9/t2/t1/p_1_in [7]),
        .I2(\r9/t2/t1/p_0_in [7]),
        .I3(\r9/t1/t0/p_1_in [7]),
        .I4(k8b[95]),
        .I5(\r9/t3/t2/p_0_in [7]),
        .O(\r9/p_0_out [95]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair343" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[95]_i_1__8 
       (.I0(\a10/k1a [31]),
        .I1(\a10/k4a [31]),
        .I2(\rf/p_2_in [31]),
        .O(\rf/p_4_out [95]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[96]_i_1 
       (.I0(\r1/t0/t0/p_1_in [0]),
        .I1(\r1/t0/t0/p_0_in [0]),
        .I2(\r1/t2/t2/p_0_in [0]),
        .I3(\r1/t1/t1/p_0_in [0]),
        .I4(k0b[96]),
        .I5(\r1/t3/t3/p_1_in [0]),
        .O(\r1/p_0_out [96]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[96]_i_1__0 
       (.I0(\r2/t0/t0/p_1_in [0]),
        .I1(\r2/t0/t0/p_0_in [0]),
        .I2(\r2/t2/t2/p_0_in [0]),
        .I3(\r2/t1/t1/p_0_in [0]),
        .I4(k1b[96]),
        .I5(\r2/t3/t3/p_1_in [0]),
        .O(\r2/p_0_out [96]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[96]_i_1__1 
       (.I0(\r3/t0/t0/p_1_in [0]),
        .I1(\r3/t0/t0/p_0_in [0]),
        .I2(\r3/t2/t2/p_0_in [0]),
        .I3(\r3/t1/t1/p_0_in [0]),
        .I4(k2b[96]),
        .I5(\r3/t3/t3/p_1_in [0]),
        .O(\r3/p_0_out [96]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[96]_i_1__2 
       (.I0(\r4/t0/t0/p_1_in [0]),
        .I1(\r4/t0/t0/p_0_in [0]),
        .I2(\r4/t2/t2/p_0_in [0]),
        .I3(\r4/t1/t1/p_0_in [0]),
        .I4(k3b[96]),
        .I5(\r4/t3/t3/p_1_in [0]),
        .O(\r4/p_0_out [96]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[96]_i_1__3 
       (.I0(\r5/t0/t0/p_1_in [0]),
        .I1(\r5/t0/t0/p_0_in [0]),
        .I2(\r5/t2/t2/p_0_in [0]),
        .I3(\r5/t1/t1/p_0_in [0]),
        .I4(k4b[96]),
        .I5(\r5/t3/t3/p_1_in [0]),
        .O(\r5/p_0_out [96]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[96]_i_1__4 
       (.I0(\r6/t0/t0/p_1_in [0]),
        .I1(\r6/t0/t0/p_0_in [0]),
        .I2(\r6/t2/t2/p_0_in [0]),
        .I3(\r6/t1/t1/p_0_in [0]),
        .I4(k5b[96]),
        .I5(\r6/t3/t3/p_1_in [0]),
        .O(\r6/p_0_out [96]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[96]_i_1__5 
       (.I0(\r7/t0/t0/p_1_in [0]),
        .I1(\r7/t0/t0/p_0_in [0]),
        .I2(\r7/t2/t2/p_0_in [0]),
        .I3(\r7/t1/t1/p_0_in [0]),
        .I4(k6b[96]),
        .I5(\r7/t3/t3/p_1_in [0]),
        .O(\r7/p_0_out [96]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[96]_i_1__6 
       (.I0(\r8/t0/t0/p_1_in [0]),
        .I1(\r8/t0/t0/p_0_in [0]),
        .I2(\r8/t2/t2/p_0_in [0]),
        .I3(\r8/t1/t1/p_0_in [0]),
        .I4(k7b[96]),
        .I5(\r8/t3/t3/p_1_in [0]),
        .O(\r8/p_0_out [96]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[96]_i_1__7 
       (.I0(\r9/t0/t0/p_1_in [0]),
        .I1(\r9/t0/t0/p_0_in [0]),
        .I2(\r9/t2/t2/p_0_in [0]),
        .I3(\r9/t1/t1/p_0_in [0]),
        .I4(k8b[96]),
        .I5(\r9/t3/t3/p_1_in [0]),
        .O(\r9/p_0_out [96]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair342" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[96]_i_1__8 
       (.I0(\a10/k0a [0]),
        .I1(\a10/k4a [0]),
        .I2(\rf/p_3_in [0]),
        .O(\rf/p_4_out [96]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[97]_i_1 
       (.I0(\r1/t0/t0/p_1_in [1]),
        .I1(\r1/t0/t0/p_0_in [1]),
        .I2(\r1/t2/t2/p_0_in [1]),
        .I3(\r1/t1/t1/p_0_in [1]),
        .I4(k0b[97]),
        .I5(\r1/t3/t3/p_1_in [1]),
        .O(\r1/p_0_out [97]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[97]_i_1__0 
       (.I0(\r2/t0/t0/p_1_in [1]),
        .I1(\r2/t0/t0/p_0_in [1]),
        .I2(\r2/t2/t2/p_0_in [1]),
        .I3(\r2/t1/t1/p_0_in [1]),
        .I4(k1b[97]),
        .I5(\r2/t3/t3/p_1_in [1]),
        .O(\r2/p_0_out [97]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[97]_i_1__1 
       (.I0(\r3/t0/t0/p_1_in [1]),
        .I1(\r3/t0/t0/p_0_in [1]),
        .I2(\r3/t2/t2/p_0_in [1]),
        .I3(\r3/t1/t1/p_0_in [1]),
        .I4(k2b[97]),
        .I5(\r3/t3/t3/p_1_in [1]),
        .O(\r3/p_0_out [97]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[97]_i_1__2 
       (.I0(\r4/t0/t0/p_1_in [1]),
        .I1(\r4/t0/t0/p_0_in [1]),
        .I2(\r4/t2/t2/p_0_in [1]),
        .I3(\r4/t1/t1/p_0_in [1]),
        .I4(k3b[97]),
        .I5(\r4/t3/t3/p_1_in [1]),
        .O(\r4/p_0_out [97]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[97]_i_1__3 
       (.I0(\r5/t0/t0/p_1_in [1]),
        .I1(\r5/t0/t0/p_0_in [1]),
        .I2(\r5/t2/t2/p_0_in [1]),
        .I3(\r5/t1/t1/p_0_in [1]),
        .I4(k4b[97]),
        .I5(\r5/t3/t3/p_1_in [1]),
        .O(\r5/p_0_out [97]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[97]_i_1__4 
       (.I0(\r6/t0/t0/p_1_in [1]),
        .I1(\r6/t0/t0/p_0_in [1]),
        .I2(\r6/t2/t2/p_0_in [1]),
        .I3(\r6/t1/t1/p_0_in [1]),
        .I4(k5b[97]),
        .I5(\r6/t3/t3/p_1_in [1]),
        .O(\r6/p_0_out [97]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[97]_i_1__5 
       (.I0(\r7/t0/t0/p_1_in [1]),
        .I1(\r7/t0/t0/p_0_in [1]),
        .I2(\r7/t2/t2/p_0_in [1]),
        .I3(\r7/t1/t1/p_0_in [1]),
        .I4(k6b[97]),
        .I5(\r7/t3/t3/p_1_in [1]),
        .O(\r7/p_0_out [97]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[97]_i_1__6 
       (.I0(\r8/t0/t0/p_1_in [1]),
        .I1(\r8/t0/t0/p_0_in [1]),
        .I2(\r8/t2/t2/p_0_in [1]),
        .I3(\r8/t1/t1/p_0_in [1]),
        .I4(k7b[97]),
        .I5(\r8/t3/t3/p_1_in [1]),
        .O(\r8/p_0_out [97]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[97]_i_1__7 
       (.I0(\r9/t0/t0/p_1_in [1]),
        .I1(\r9/t0/t0/p_0_in [1]),
        .I2(\r9/t2/t2/p_0_in [1]),
        .I3(\r9/t1/t1/p_0_in [1]),
        .I4(k8b[97]),
        .I5(\r9/t3/t3/p_1_in [1]),
        .O(\r9/p_0_out [97]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair341" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[97]_i_1__8 
       (.I0(\a10/k0a [1]),
        .I1(\a10/k4a [1]),
        .I2(\rf/p_3_in [1]),
        .O(\rf/p_4_out [97]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[98]_i_1 
       (.I0(\r1/t0/t0/p_1_in [2]),
        .I1(\r1/t0/t0/p_0_in [2]),
        .I2(\r1/t2/t2/p_0_in [2]),
        .I3(\r1/t1/t1/p_0_in [2]),
        .I4(k0b[98]),
        .I5(\r1/t3/t3/p_1_in [2]),
        .O(\r1/p_0_out [98]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[98]_i_1__0 
       (.I0(\r2/t0/t0/p_1_in [2]),
        .I1(\r2/t0/t0/p_0_in [2]),
        .I2(\r2/t2/t2/p_0_in [2]),
        .I3(\r2/t1/t1/p_0_in [2]),
        .I4(k1b[98]),
        .I5(\r2/t3/t3/p_1_in [2]),
        .O(\r2/p_0_out [98]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[98]_i_1__1 
       (.I0(\r3/t0/t0/p_1_in [2]),
        .I1(\r3/t0/t0/p_0_in [2]),
        .I2(\r3/t2/t2/p_0_in [2]),
        .I3(\r3/t1/t1/p_0_in [2]),
        .I4(k2b[98]),
        .I5(\r3/t3/t3/p_1_in [2]),
        .O(\r3/p_0_out [98]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[98]_i_1__2 
       (.I0(\r4/t0/t0/p_1_in [2]),
        .I1(\r4/t0/t0/p_0_in [2]),
        .I2(\r4/t2/t2/p_0_in [2]),
        .I3(\r4/t1/t1/p_0_in [2]),
        .I4(k3b[98]),
        .I5(\r4/t3/t3/p_1_in [2]),
        .O(\r4/p_0_out [98]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[98]_i_1__3 
       (.I0(\r5/t0/t0/p_1_in [2]),
        .I1(\r5/t0/t0/p_0_in [2]),
        .I2(\r5/t2/t2/p_0_in [2]),
        .I3(\r5/t1/t1/p_0_in [2]),
        .I4(k4b[98]),
        .I5(\r5/t3/t3/p_1_in [2]),
        .O(\r5/p_0_out [98]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[98]_i_1__4 
       (.I0(\r6/t0/t0/p_1_in [2]),
        .I1(\r6/t0/t0/p_0_in [2]),
        .I2(\r6/t2/t2/p_0_in [2]),
        .I3(\r6/t1/t1/p_0_in [2]),
        .I4(k5b[98]),
        .I5(\r6/t3/t3/p_1_in [2]),
        .O(\r6/p_0_out [98]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[98]_i_1__5 
       (.I0(\r7/t0/t0/p_1_in [2]),
        .I1(\r7/t0/t0/p_0_in [2]),
        .I2(\r7/t2/t2/p_0_in [2]),
        .I3(\r7/t1/t1/p_0_in [2]),
        .I4(k6b[98]),
        .I5(\r7/t3/t3/p_1_in [2]),
        .O(\r7/p_0_out [98]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[98]_i_1__6 
       (.I0(\r8/t0/t0/p_1_in [2]),
        .I1(\r8/t0/t0/p_0_in [2]),
        .I2(\r8/t2/t2/p_0_in [2]),
        .I3(\r8/t1/t1/p_0_in [2]),
        .I4(k7b[98]),
        .I5(\r8/t3/t3/p_1_in [2]),
        .O(\r8/p_0_out [98]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[98]_i_1__7 
       (.I0(\r9/t0/t0/p_1_in [2]),
        .I1(\r9/t0/t0/p_0_in [2]),
        .I2(\r9/t2/t2/p_0_in [2]),
        .I3(\r9/t1/t1/p_0_in [2]),
        .I4(k8b[98]),
        .I5(\r9/t3/t3/p_1_in [2]),
        .O(\r9/p_0_out [98]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair340" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[98]_i_1__8 
       (.I0(\a10/k0a [2]),
        .I1(\a10/k4a [2]),
        .I2(\rf/p_3_in [2]),
        .O(\rf/p_4_out [98]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[99]_i_1 
       (.I0(\r1/t0/t0/p_1_in [3]),
        .I1(\r1/t0/t0/p_0_in [3]),
        .I2(\r1/t2/t2/p_0_in [3]),
        .I3(\r1/t1/t1/p_0_in [3]),
        .I4(k0b[99]),
        .I5(\r1/t3/t3/p_1_in [3]),
        .O(\r1/p_0_out [99]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[99]_i_1__0 
       (.I0(\r2/t0/t0/p_1_in [3]),
        .I1(\r2/t0/t0/p_0_in [3]),
        .I2(\r2/t2/t2/p_0_in [3]),
        .I3(\r2/t1/t1/p_0_in [3]),
        .I4(k1b[99]),
        .I5(\r2/t3/t3/p_1_in [3]),
        .O(\r2/p_0_out [99]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[99]_i_1__1 
       (.I0(\r3/t0/t0/p_1_in [3]),
        .I1(\r3/t0/t0/p_0_in [3]),
        .I2(\r3/t2/t2/p_0_in [3]),
        .I3(\r3/t1/t1/p_0_in [3]),
        .I4(k2b[99]),
        .I5(\r3/t3/t3/p_1_in [3]),
        .O(\r3/p_0_out [99]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[99]_i_1__2 
       (.I0(\r4/t0/t0/p_1_in [3]),
        .I1(\r4/t0/t0/p_0_in [3]),
        .I2(\r4/t2/t2/p_0_in [3]),
        .I3(\r4/t1/t1/p_0_in [3]),
        .I4(k3b[99]),
        .I5(\r4/t3/t3/p_1_in [3]),
        .O(\r4/p_0_out [99]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[99]_i_1__3 
       (.I0(\r5/t0/t0/p_1_in [3]),
        .I1(\r5/t0/t0/p_0_in [3]),
        .I2(\r5/t2/t2/p_0_in [3]),
        .I3(\r5/t1/t1/p_0_in [3]),
        .I4(k4b[99]),
        .I5(\r5/t3/t3/p_1_in [3]),
        .O(\r5/p_0_out [99]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[99]_i_1__4 
       (.I0(\r6/t0/t0/p_1_in [3]),
        .I1(\r6/t0/t0/p_0_in [3]),
        .I2(\r6/t2/t2/p_0_in [3]),
        .I3(\r6/t1/t1/p_0_in [3]),
        .I4(k5b[99]),
        .I5(\r6/t3/t3/p_1_in [3]),
        .O(\r6/p_0_out [99]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[99]_i_1__5 
       (.I0(\r7/t0/t0/p_1_in [3]),
        .I1(\r7/t0/t0/p_0_in [3]),
        .I2(\r7/t2/t2/p_0_in [3]),
        .I3(\r7/t1/t1/p_0_in [3]),
        .I4(k6b[99]),
        .I5(\r7/t3/t3/p_1_in [3]),
        .O(\r7/p_0_out [99]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[99]_i_1__6 
       (.I0(\r8/t0/t0/p_1_in [3]),
        .I1(\r8/t0/t0/p_0_in [3]),
        .I2(\r8/t2/t2/p_0_in [3]),
        .I3(\r8/t1/t1/p_0_in [3]),
        .I4(k7b[99]),
        .I5(\r8/t3/t3/p_1_in [3]),
        .O(\r8/p_0_out [99]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[99]_i_1__7 
       (.I0(\r9/t0/t0/p_1_in [3]),
        .I1(\r9/t0/t0/p_0_in [3]),
        .I2(\r9/t2/t2/p_0_in [3]),
        .I3(\r9/t1/t1/p_0_in [3]),
        .I4(k8b[99]),
        .I5(\r9/t3/t3/p_1_in [3]),
        .O(\r9/p_0_out [99]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair339" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[99]_i_1__8 
       (.I0(\a10/k0a [3]),
        .I1(\a10/k4a [3]),
        .I2(\rf/p_3_in [3]),
        .O(\rf/p_4_out [99]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[9]_i_1 
       (.I0(\r1/t0/t1/p_0_in [1]),
        .I1(\r1/t2/t3/p_1_in [1]),
        .I2(\r1/t2/t3/p_0_in [1]),
        .I3(\r1/t1/t2/p_1_in [1]),
        .I4(k0b[9]),
        .I5(\r1/t3/t0/p_0_in [1]),
        .O(\r1/p_0_out [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[9]_i_1__0 
       (.I0(\r2/t0/t1/p_0_in [1]),
        .I1(\r2/t2/t3/p_1_in [1]),
        .I2(\r2/t2/t3/p_0_in [1]),
        .I3(\r2/t1/t2/p_1_in [1]),
        .I4(k1b[9]),
        .I5(\r2/t3/t0/p_0_in [1]),
        .O(\r2/p_0_out [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[9]_i_1__1 
       (.I0(\r3/t0/t1/p_0_in [1]),
        .I1(\r3/t2/t3/p_1_in [1]),
        .I2(\r3/t2/t3/p_0_in [1]),
        .I3(\r3/t1/t2/p_1_in [1]),
        .I4(k2b[9]),
        .I5(\r3/t3/t0/p_0_in [1]),
        .O(\r3/p_0_out [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[9]_i_1__2 
       (.I0(\r4/t0/t1/p_0_in [1]),
        .I1(\r4/t2/t3/p_1_in [1]),
        .I2(\r4/t2/t3/p_0_in [1]),
        .I3(\r4/t1/t2/p_1_in [1]),
        .I4(k3b[9]),
        .I5(\r4/t3/t0/p_0_in [1]),
        .O(\r4/p_0_out [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[9]_i_1__3 
       (.I0(\r5/t0/t1/p_0_in [1]),
        .I1(\r5/t2/t3/p_1_in [1]),
        .I2(\r5/t2/t3/p_0_in [1]),
        .I3(\r5/t1/t2/p_1_in [1]),
        .I4(k4b[9]),
        .I5(\r5/t3/t0/p_0_in [1]),
        .O(\r5/p_0_out [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[9]_i_1__4 
       (.I0(\r6/t0/t1/p_0_in [1]),
        .I1(\r6/t2/t3/p_1_in [1]),
        .I2(\r6/t2/t3/p_0_in [1]),
        .I3(\r6/t1/t2/p_1_in [1]),
        .I4(k5b[9]),
        .I5(\r6/t3/t0/p_0_in [1]),
        .O(\r6/p_0_out [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[9]_i_1__5 
       (.I0(\r7/t0/t1/p_0_in [1]),
        .I1(\r7/t2/t3/p_1_in [1]),
        .I2(\r7/t2/t3/p_0_in [1]),
        .I3(\r7/t1/t2/p_1_in [1]),
        .I4(k6b[9]),
        .I5(\r7/t3/t0/p_0_in [1]),
        .O(\r7/p_0_out [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[9]_i_1__6 
       (.I0(\r8/t0/t1/p_0_in [1]),
        .I1(\r8/t2/t3/p_1_in [1]),
        .I2(\r8/t2/t3/p_0_in [1]),
        .I3(\r8/t1/t2/p_1_in [1]),
        .I4(k7b[9]),
        .I5(\r8/t3/t0/p_0_in [1]),
        .O(\r8/p_0_out [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \state_out[9]_i_1__7 
       (.I0(\r9/t0/t1/p_0_in [1]),
        .I1(\r9/t2/t3/p_1_in [1]),
        .I2(\r9/t2/t3/p_0_in [1]),
        .I3(\r9/t1/t2/p_1_in [1]),
        .I4(k8b[9]),
        .I5(\r9/t3/t0/p_0_in [1]),
        .O(\r9/p_0_out [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair333" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \state_out[9]_i_1__8 
       (.I0(\a10/k3a [9]),
        .I1(\a10/k4a [9]),
        .I2(\rf/p_0_in [9]),
        .O(\rf/p_4_out [9]));
endmodule
