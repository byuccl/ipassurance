module fixed_point_sqrt
   (clk,
    res,
    ARG,
    backdoor,
    Z);
  output backdoor;
  input clk;
  input res;
  input [31:0]ARG;
  output [31:0]Z;

  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const0>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const1>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]ARG;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire GND_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire RSTA;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire VCC_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]Z;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire clk;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\d_next[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [47:0]d_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_106 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_107 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_108 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_109 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_111 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_112 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_113 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_114 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_115 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_116 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_117 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_118 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_119 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_121 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_122 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_123 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_124 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_125 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_126 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_127 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_128 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_129 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_131 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_132 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_133 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_134 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_135 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_136 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_137 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_138 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_139 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_141 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_142 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_143 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_144 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_145 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_146 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_147 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_148 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_149 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_150 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_151 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_152 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_153 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__1_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__2_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0__2_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_10__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_11__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_12__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_13__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_14__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_6__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_7__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_8__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_9__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_106 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_107 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_108 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_109 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_111 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_112 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_113 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_114 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_115 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_116 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_117 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_118 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_119 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_121 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_122 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_123 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_124 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_125 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_126 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_127 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_128 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_129 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_131 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_132 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_133 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_134 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_135 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_136 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_137 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_138 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_139 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_141 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_142 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_143 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_144 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_145 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_146 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_147 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_148 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_149 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_150 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_151 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_152 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_153 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \d_reg[1]0_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b10__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b11__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b12__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b13__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b14__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b15__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b16__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b17__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b18__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b19__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b20__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b21__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b22__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b23__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b24__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b24_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b25__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b25_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b26__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b26_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b27__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b27_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b28__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b28_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b29__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b29_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b30_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b5__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b6__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b7__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b8__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b9__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b0__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b10__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b11__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b12__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b13__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b14__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b15__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b16__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b17__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b18__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b19__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b20__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b21__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b22__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b23__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b24__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b24_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b25__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b25_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b26__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b26_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b27__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b27_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b28__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b28_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b29_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b5__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b6__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b7__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b8__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b9__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire n;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][0]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][0]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][0]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][0]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][0]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][0]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][0]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][0]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][16]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][16]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][16]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][16]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][20]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][20]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][20]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][20]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][24]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][24]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][24]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][24]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][28]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][28]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][28]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][28]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][31]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n[3][8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\n_next[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\n_next[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\n_next[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [47:0]n_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_106 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_107 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_108 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_109 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_111 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_112 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_113 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_114 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_115 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_116 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_117 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_118 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_119 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_121 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_122 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_123 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_124 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_125 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_126 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_127 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_128 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_129 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_131 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_132 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_133 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_134 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_135 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_136 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_137 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_138 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_139 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_141 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_142 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_143 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_144 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_145 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_146 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_147 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_148 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_149 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_150 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_151 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_152 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_153 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__1_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0__2_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_10__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_11__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_12__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_6__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_7__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_8__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_9__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_106 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_107 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_108 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_109 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_111 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_112 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_113 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_114 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_115 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_116 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_117 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_118 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_119 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_121 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_122 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_123 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_124 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_125 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_126 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_127 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_128 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_129 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_131 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_132 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_133 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_134 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_135 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_136 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_137 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_138 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_139 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_141 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_142 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_143 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_144 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_145 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_146 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_147 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_148 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_149 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_150 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_151 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_152 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_153 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[1]0_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__0_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_106 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_107 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_108 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_109 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_111 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_112 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_113 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_114 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_115 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_116 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_117 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_118 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_119 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_121 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_122 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_123 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_124 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_125 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_126 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_127 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_128 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_129 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_131 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_132 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_133 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_134 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_135 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_136 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_137 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_138 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_139 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_141 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_142 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_143 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_144 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_145 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_146 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_147 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_148 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_149 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_150 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_151 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_152 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_153 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_24 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_25 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_26 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_27 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_28 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_29 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_30 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_31 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_32 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_33 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_34 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_35 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_36 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_37 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_38 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_39 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_40 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_41 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_42 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_43 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_44 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_45 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_46 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_47 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_48 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_49 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_50 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_51 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_52 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_53 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__1_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0__2_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_10__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_11__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_12__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_13__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_14__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_15__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_16__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_17__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_18__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_19__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_1__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_22_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_22_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_22_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_27_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_27_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_27_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_2__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_2__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_2__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_32_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_32_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_3__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_3__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_3__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_4__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_4__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_4__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_4_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_5_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_5_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_5_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_5_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_5_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_5_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_6__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_7__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_8__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_9__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_106 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_107 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_108 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_109 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_111 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_112 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_113 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_114 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_115 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_116 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_117 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_118 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_119 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_121 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_122 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_123 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_124 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_125 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_126 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_127 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_128 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_129 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_131 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_132 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_133 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_134 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_135 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_136 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_137 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_138 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_139 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_141 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_142 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_143 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_144 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_145 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_146 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_147 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_148 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_149 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_150 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_151 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_152 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_153 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[2]0_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__0_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_106 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_107 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_108 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_109 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_111 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_112 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_113 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_114 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_115 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_116 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_117 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_118 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_119 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_121 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_122 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_123 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_124 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_125 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_126 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_127 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_128 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_129 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_131 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_132 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_133 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_134 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_135 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_136 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_137 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_138 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_139 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_141 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_142 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_143 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_144 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_145 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_146 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_147 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_148 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_149 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_150 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_151 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_152 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_153 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_24 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_25 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_26 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_27 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_28 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_29 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_30 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_31 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_32 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_33 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_34 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_35 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_36 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_37 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_38 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_39 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_40 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_41 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_42 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_43 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_44 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_45 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_46 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_47 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_48 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_49 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_50 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_51 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_52 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_53 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__1_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0__2_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_10__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_10__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_11__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_11__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_12__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_12__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_13__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_13__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_14__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_14__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_15__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_15__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_16__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_16__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_17__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_17__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_18__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_18__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_19__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_19__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_1__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_1__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_1__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_1__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_1__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_20__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_20__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_20__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_20__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_20__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_21__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_21__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_21__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_21__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_21__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_21__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_21__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_21__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_21__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_22__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_22__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_22__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_22__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_22__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_22__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_22__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_22__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_22__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_22_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_22_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_22_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_23__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_23__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_24__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_24__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_25__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_25__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_26__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_26__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_27__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_27__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_27_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_27_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_27_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_28__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_28__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_29__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_29__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_2__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_2__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_2__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_2__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_2__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_2__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_30__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_30__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_31__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_31__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_32__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_32__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_32_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_32_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_33__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_33__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_34__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_35__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_36__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_37__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_38__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_39__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_3__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_3__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_3__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_3__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_3__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_3__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_42_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_42_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_42_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_47_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_47_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_47_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_47_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_47_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_47_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_47_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_48_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_48_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_48_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_48_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_48_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_48_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_48_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_49_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_49_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_49_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_49_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_49_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_49_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_49_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_4__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_4__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_4__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_4__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_4__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_4__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_4__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_4_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_50_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_50_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_50_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_50_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_50_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_50_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_50_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_51_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_51_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_51_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_52_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_53_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_54_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_55_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_57_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_58_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_59_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_5__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_5__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_5__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_5__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_5_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_5_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_5_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_5_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_5_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_5_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_60_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_61_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_62_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_63_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_64_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_65_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_66_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_67_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_68_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_69_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_6__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_6__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_6__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_6__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_70_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_71_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_72_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_72_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_72_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_72_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_73_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_74_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_75_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_76_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_77_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_77_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_77_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_77_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_78_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_79_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_7__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_7__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_7__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_7__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_7__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_80_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_81_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_82_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_83_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_84_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_8__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_8__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_8__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_8__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_8__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_9__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_9__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_9__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_9__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_9__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_9__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_9__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_9__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_9__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_106 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_107 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_108 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_109 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_111 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_112 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_113 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_114 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_115 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_116 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_117 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_118 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_119 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_121 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_122 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_123 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_124 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_125 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_126 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_127 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_128 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_129 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_131 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_132 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_133 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_134 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_135 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_136 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_137 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_138 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_139 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_141 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_142 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_143 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_144 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_145 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_146 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_147 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_148 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_149 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_150 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_151 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_152 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_153 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3]0_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][0]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][0]_i_12_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][0]_i_12_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][0]_i_12_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][0]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][0]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][0]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][0]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][0]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][0]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][0]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][0]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][0]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][0]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][0]_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][0]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][12]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][12]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][12]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][16]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][16]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][16]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][20]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][20]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][20]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][24]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][24]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][24]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][28]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][28]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][28]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][31]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][4]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][4]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][4]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][8]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][8]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \n_reg[3][8]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [30:0]p_0_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [62:16]p_1_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_10;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_11;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_12;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_13;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_14;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_15;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_16;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_17;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_18;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_19;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_20;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_21;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_22;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_23;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_24;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_25;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_26;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_27;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_28;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_29;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_30;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_31;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_32;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_33;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_34;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_35;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_36;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_37;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_38;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_39;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_4;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_40;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_41;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_42;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_43;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_44;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_45;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_46;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_47;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_48;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_49;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_5;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_50;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_51;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_52;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_53;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_54;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_55;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_56;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_57;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_58;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_59;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_6;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_60;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_61;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_62;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_63;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_7;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_8;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire psdsp_n_9;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [47:0]r_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:1]\r_reg[1]0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:1]\r_reg[2]0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_106 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_107 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_108 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_109 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_111 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_112 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_113 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_114 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_115 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_116 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_117 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_118 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_119 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_121 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_122 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_123 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_124 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_125 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_126 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_127 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_128 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_129 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_131 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_132 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_133 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_134 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_135 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_136 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_137 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_138 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_139 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_141 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_142 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_143 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_144 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_145 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_146 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_147 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_148 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_149 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_150 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_151 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_152 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_153 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__1_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1__2_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_10__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_10__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_11__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_11__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_12__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_12__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_13__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_13__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_14__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_14__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_15__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_15__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_16__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_16__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_17__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_17__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_17__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_17__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_17__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_18__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_18__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_19__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_19__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_1__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_1__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_1__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_1__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_20__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_21__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_22__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_22_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_22_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_22_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_23__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_24__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_25__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_26__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_27__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_27__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_27__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_27__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_28__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_29__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_2__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_2__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_2__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_2__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_2__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_2__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_30__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_31__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_32__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_33__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_34__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_3__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_3__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_3__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_3__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_3__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_3__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_41_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_41_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_41_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_46_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_46_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_46_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_4__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_4__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_4__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_4__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_4__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_4__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_4__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_4__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_4__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_4__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_4_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_51_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_51_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_51_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_52_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_53_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_54_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_55_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_57_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_58_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_5__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_5_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_5_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_5_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_6__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_6__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_6_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_6_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_6_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_7__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_7__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_8__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_8__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_8_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_8_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_9__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_9__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_9_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_9_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_9_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_9_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_9_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_i_9_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_106 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_107 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_108 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_109 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_111 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_112 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_113 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_114 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_115 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_116 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_117 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_118 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_119 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_121 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_122 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_123 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_124 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_125 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_126 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_127 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_128 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_129 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_131 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_132 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_133 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_134 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_135 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_136 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_137 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_138 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_139 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_141 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_142 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_143 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_144 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_145 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_146 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_147 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_148 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_149 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_150 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_151 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_152 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_153 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[2]1_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire res;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\rsqr_next[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [47:0]rsqr_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_106 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_107 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_108 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_109 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_111 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_112 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_113 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_114 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_115 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_116 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_117 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_118 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_119 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_121 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_122 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_123 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_124 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_125 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_126 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_127 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_128 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_129 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_131 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_132 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_133 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_134 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_135 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_136 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_137 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_138 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_139 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_141 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_142 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_143 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_144 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_145 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_146 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_147 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_148 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_149 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_150 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_151 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_152 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_153 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__1_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0__2_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_4_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_5_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_5_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_5_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_6_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_6_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_6_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_8_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_8_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_9_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_9_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_i_9_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_106 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_107 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_108 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_109 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_111 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_112 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_113 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_114 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_115 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_116 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_117 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_118 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_119 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_121 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_122 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_123 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_124 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_125 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_126 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_127 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_128 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_129 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_131 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_132 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_133 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_134 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_135 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_136 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_137 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_138 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_139 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_141 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_142 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_143 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_144 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_145 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_146 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_147 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_148 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_149 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_150 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_151 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_152 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_153 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rsqr_reg[1]0_n_99 ;

  assign backdoor =  res ;

  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND
       (.G(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_1
       (.G(GND_2));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC
       (.P(\<const1>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC_1
       (.P(VCC_2));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-10 {cell *THIS*} {string 16x18 4}}" *) 
  DSP48E1 #(
    .ACASCREG(1),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(1),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(1),
    .BREG(1),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \d_reg[1]0 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\d_reg[1]0_i_1_n_0 ,\d_reg[1]0_i_2_n_0 ,\d_reg[1]0_i_3_n_0 ,\d_reg[1]0_i_4_n_0 ,\d_reg[1]0_i_5_n_0 ,\d_reg[1]0_i_6_n_0 ,\d_reg[1]0_i_7_n_0 ,\d_reg[1]0_i_8_n_0 ,\d_reg[1]0_i_9_n_0 ,\d_reg[1]0_i_10_n_0 ,\d_reg[1]0_i_11_n_0 ,\d_reg[1]0_i_12_n_0 ,\d_reg[1]0_i_13_n_0 ,\d_reg[1]0_i_14_n_0 ,\d_reg[1]0_i_15_n_0 ,\d_reg[1]0_i_16_n_0 ,\d_reg[1]0_i_17_n_0 }),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,ARG[31:17]}),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const1>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const1>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\d_reg[1]0_n_58 ,\d_reg[1]0_n_59 ,\d_reg[1]0_n_60 ,\d_reg[1]0_n_61 ,\d_reg[1]0_n_62 ,\d_reg[1]0_n_63 ,\d_reg[1]0_n_64 ,\d_reg[1]0_n_65 ,\d_reg[1]0_n_66 ,\d_reg[1]0_n_67 ,\d_reg[1]0_n_68 ,\d_reg[1]0_n_69 ,\d_reg[1]0_n_70 ,\d_reg[1]0_n_71 ,\d_reg[1]0_n_72 ,\d_reg[1]0_n_73 ,\d_reg[1]0_n_74 ,\d_reg[1]0_n_75 ,\d_reg[1]0_n_76 ,\d_reg[1]0_n_77 ,\d_reg[1]0_n_78 ,\d_reg[1]0_n_79 ,\d_reg[1]0_n_80 ,\d_reg[1]0_n_81 ,\d_reg[1]0_n_82 ,\d_reg[1]0_n_83 ,\d_reg[1]0_n_84 ,\d_reg[1]0_n_85 ,\d_reg[1]0_n_86 ,\d_reg[1]0_n_87 ,\d_reg[1]0_n_88 ,\d_reg[1]0_n_89 ,\d_reg[1]0_n_90 ,\d_reg[1]0_n_91 ,\d_reg[1]0_n_92 ,\d_reg[1]0_n_93 ,\d_reg[1]0_n_94 ,\d_reg[1]0_n_95 ,\d_reg[1]0_n_96 ,\d_reg[1]0_n_97 ,\d_reg[1]0_n_98 ,\d_reg[1]0_n_99 ,\d_reg[1]0_n_100 ,\d_reg[1]0_n_101 ,\d_reg[1]0_n_102 ,\d_reg[1]0_n_103 ,\d_reg[1]0_n_104 ,\d_reg[1]0_n_105 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .PCOUT({\d_reg[1]0_n_106 ,\d_reg[1]0_n_107 ,\d_reg[1]0_n_108 ,\d_reg[1]0_n_109 ,\d_reg[1]0_n_110 ,\d_reg[1]0_n_111 ,\d_reg[1]0_n_112 ,\d_reg[1]0_n_113 ,\d_reg[1]0_n_114 ,\d_reg[1]0_n_115 ,\d_reg[1]0_n_116 ,\d_reg[1]0_n_117 ,\d_reg[1]0_n_118 ,\d_reg[1]0_n_119 ,\d_reg[1]0_n_120 ,\d_reg[1]0_n_121 ,\d_reg[1]0_n_122 ,\d_reg[1]0_n_123 ,\d_reg[1]0_n_124 ,\d_reg[1]0_n_125 ,\d_reg[1]0_n_126 ,\d_reg[1]0_n_127 ,\d_reg[1]0_n_128 ,\d_reg[1]0_n_129 ,\d_reg[1]0_n_130 ,\d_reg[1]0_n_131 ,\d_reg[1]0_n_132 ,\d_reg[1]0_n_133 ,\d_reg[1]0_n_134 ,\d_reg[1]0_n_135 ,\d_reg[1]0_n_136 ,\d_reg[1]0_n_137 ,\d_reg[1]0_n_138 ,\d_reg[1]0_n_139 ,\d_reg[1]0_n_140 ,\d_reg[1]0_n_141 ,\d_reg[1]0_n_142 ,\d_reg[1]0_n_143 ,\d_reg[1]0_n_144 ,\d_reg[1]0_n_145 ,\d_reg[1]0_n_146 ,\d_reg[1]0_n_147 ,\d_reg[1]0_n_148 ,\d_reg[1]0_n_149 ,\d_reg[1]0_n_150 ,\d_reg[1]0_n_151 ,\d_reg[1]0_n_152 ,\d_reg[1]0_n_153 }),
        .RSTA(RSTA),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(RSTA),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-10 {cell *THIS*} {string 16x16 4}}" *) 
  DSP48E1 #(
    .ACASCREG(1),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(1),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(1),
    .BREG(1),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \d_reg[1]0__0 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,ARG[31:17]}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\d_reg[1]0_i_1__0_n_0 ,\d_reg[1]0_i_2__0_n_0 ,\d_reg[1]0_i_3__0_n_0 ,\d_reg[1]0_i_4__0_n_0 ,\d_reg[1]0_i_5__0_n_0 ,\d_reg[1]0_i_6__0_n_0 ,\d_reg[1]0_i_7__0_n_0 ,\d_reg[1]0_i_8__0_n_0 ,\d_reg[1]0_i_9__0_n_0 ,\d_reg[1]0_i_10__0_n_0 ,\d_reg[1]0_i_11__0_n_0 ,\d_reg[1]0_i_12__0_n_0 ,\d_reg[1]0_i_13__0_n_0 ,\d_reg[1]0_i_14__0_n_0 }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const1>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const1>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P(d_reg),
        .PCIN({\d_reg[1]0_n_106 ,\d_reg[1]0_n_107 ,\d_reg[1]0_n_108 ,\d_reg[1]0_n_109 ,\d_reg[1]0_n_110 ,\d_reg[1]0_n_111 ,\d_reg[1]0_n_112 ,\d_reg[1]0_n_113 ,\d_reg[1]0_n_114 ,\d_reg[1]0_n_115 ,\d_reg[1]0_n_116 ,\d_reg[1]0_n_117 ,\d_reg[1]0_n_118 ,\d_reg[1]0_n_119 ,\d_reg[1]0_n_120 ,\d_reg[1]0_n_121 ,\d_reg[1]0_n_122 ,\d_reg[1]0_n_123 ,\d_reg[1]0_n_124 ,\d_reg[1]0_n_125 ,\d_reg[1]0_n_126 ,\d_reg[1]0_n_127 ,\d_reg[1]0_n_128 ,\d_reg[1]0_n_129 ,\d_reg[1]0_n_130 ,\d_reg[1]0_n_131 ,\d_reg[1]0_n_132 ,\d_reg[1]0_n_133 ,\d_reg[1]0_n_134 ,\d_reg[1]0_n_135 ,\d_reg[1]0_n_136 ,\d_reg[1]0_n_137 ,\d_reg[1]0_n_138 ,\d_reg[1]0_n_139 ,\d_reg[1]0_n_140 ,\d_reg[1]0_n_141 ,\d_reg[1]0_n_142 ,\d_reg[1]0_n_143 ,\d_reg[1]0_n_144 ,\d_reg[1]0_n_145 ,\d_reg[1]0_n_146 ,\d_reg[1]0_n_147 ,\d_reg[1]0_n_148 ,\d_reg[1]0_n_149 ,\d_reg[1]0_n_150 ,\d_reg[1]0_n_151 ,\d_reg[1]0_n_152 ,\d_reg[1]0_n_153 }),
        .RSTA(RSTA),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(RSTA),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-10 {cell *THIS*} {string 18x18 4}}" *) 
  DSP48E1 #(
    .ACASCREG(1),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(1),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(1),
    .BREG(1),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \d_reg[1]0__1 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,ARG[16:0]}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\d_reg[1]0_i_1_n_0 ,\d_reg[1]0_i_2_n_0 ,\d_reg[1]0_i_3_n_0 ,\d_reg[1]0_i_4_n_0 ,\d_reg[1]0_i_5_n_0 ,\d_reg[1]0_i_6_n_0 ,\d_reg[1]0_i_7_n_0 ,\d_reg[1]0_i_8_n_0 ,\d_reg[1]0_i_9_n_0 ,\d_reg[1]0_i_10_n_0 ,\d_reg[1]0_i_11_n_0 ,\d_reg[1]0_i_12_n_0 ,\d_reg[1]0_i_13_n_0 ,\d_reg[1]0_i_14_n_0 ,\d_reg[1]0_i_15_n_0 ,\d_reg[1]0_i_16_n_0 ,\d_reg[1]0_i_17_n_0 }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const1>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const1>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\d_reg[1]0__1_n_58 ,\d_reg[1]0__1_n_59 ,\d_reg[1]0__1_n_60 ,\d_reg[1]0__1_n_61 ,\d_reg[1]0__1_n_62 ,\d_reg[1]0__1_n_63 ,\d_reg[1]0__1_n_64 ,\d_reg[1]0__1_n_65 ,\d_reg[1]0__1_n_66 ,\d_reg[1]0__1_n_67 ,\d_reg[1]0__1_n_68 ,\d_reg[1]0__1_n_69 ,\d_reg[1]0__1_n_70 ,\d_reg[1]0__1_n_71 ,\d_reg[1]0__1_n_72 ,\d_reg[1]0__1_n_73 ,\d_reg[1]0__1_n_74 ,\d_reg[1]0__1_n_75 ,\d_reg[1]0__1_n_76 ,\d_reg[1]0__1_n_77 ,\d_reg[1]0__1_n_78 ,\d_reg[1]0__1_n_79 ,\d_reg[1]0__1_n_80 ,\d_reg[1]0__1_n_81 ,\d_reg[1]0__1_n_82 ,\d_reg[1]0__1_n_83 ,\d_reg[1]0__1_n_84 ,\d_reg[1]0__1_n_85 ,\d_reg[1]0__1_n_86 ,\d_reg[1]0__1_n_87 ,\d_reg[1]0__1_n_88 ,p_1_in[16],\d_reg[1]0__1_n_90 ,\d_reg[1]0__1_n_91 ,\d_reg[1]0__1_n_92 ,\d_reg[1]0__1_n_93 ,\d_reg[1]0__1_n_94 ,\d_reg[1]0__1_n_95 ,\d_reg[1]0__1_n_96 ,\d_reg[1]0__1_n_97 ,\d_reg[1]0__1_n_98 ,\d_reg[1]0__1_n_99 ,\d_reg[1]0__1_n_100 ,\d_reg[1]0__1_n_101 ,\d_reg[1]0__1_n_102 ,\d_reg[1]0__1_n_103 ,\d_reg[1]0__1_n_104 ,\d_reg[1]0__1_n_105 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .PCOUT({\d_reg[1]0__1_n_106 ,\d_reg[1]0__1_n_107 ,\d_reg[1]0__1_n_108 ,\d_reg[1]0__1_n_109 ,\d_reg[1]0__1_n_110 ,\d_reg[1]0__1_n_111 ,\d_reg[1]0__1_n_112 ,\d_reg[1]0__1_n_113 ,\d_reg[1]0__1_n_114 ,\d_reg[1]0__1_n_115 ,\d_reg[1]0__1_n_116 ,\d_reg[1]0__1_n_117 ,\d_reg[1]0__1_n_118 ,\d_reg[1]0__1_n_119 ,\d_reg[1]0__1_n_120 ,\d_reg[1]0__1_n_121 ,\d_reg[1]0__1_n_122 ,\d_reg[1]0__1_n_123 ,\d_reg[1]0__1_n_124 ,\d_reg[1]0__1_n_125 ,\d_reg[1]0__1_n_126 ,\d_reg[1]0__1_n_127 ,\d_reg[1]0__1_n_128 ,\d_reg[1]0__1_n_129 ,\d_reg[1]0__1_n_130 ,\d_reg[1]0__1_n_131 ,\d_reg[1]0__1_n_132 ,\d_reg[1]0__1_n_133 ,\d_reg[1]0__1_n_134 ,\d_reg[1]0__1_n_135 ,\d_reg[1]0__1_n_136 ,\d_reg[1]0__1_n_137 ,\d_reg[1]0__1_n_138 ,\d_reg[1]0__1_n_139 ,\d_reg[1]0__1_n_140 ,\d_reg[1]0__1_n_141 ,\d_reg[1]0__1_n_142 ,\d_reg[1]0__1_n_143 ,\d_reg[1]0__1_n_144 ,\d_reg[1]0__1_n_145 ,\d_reg[1]0__1_n_146 ,\d_reg[1]0__1_n_147 ,\d_reg[1]0__1_n_148 ,\d_reg[1]0__1_n_149 ,\d_reg[1]0__1_n_150 ,\d_reg[1]0__1_n_151 ,\d_reg[1]0__1_n_152 ,\d_reg[1]0__1_n_153 }),
        .RSTA(RSTA),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(RSTA),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-10 {cell *THIS*} {string 18x16 4}}" *) 
  DSP48E1 #(
    .ACASCREG(1),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(1),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(1),
    .BREG(1),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \d_reg[1]0__2 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,ARG[16:0]}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\d_reg[1]0_i_1__0_n_0 ,\d_reg[1]0_i_2__0_n_0 ,\d_reg[1]0_i_3__0_n_0 ,\d_reg[1]0_i_4__0_n_0 ,\d_reg[1]0_i_5__0_n_0 ,\d_reg[1]0_i_6__0_n_0 ,\d_reg[1]0_i_7__0_n_0 ,\d_reg[1]0_i_8__0_n_0 ,\d_reg[1]0_i_9__0_n_0 ,\d_reg[1]0_i_10__0_n_0 ,\d_reg[1]0_i_11__0_n_0 ,\d_reg[1]0_i_12__0_n_0 ,\d_reg[1]0_i_13__0_n_0 ,\d_reg[1]0_i_14__0_n_0 }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const1>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const1>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\d_reg[1]0__2_n_58 ,\d_reg[1]0__2_n_59 ,p_1_in[62:17]}),
        .PCIN({\d_reg[1]0__1_n_106 ,\d_reg[1]0__1_n_107 ,\d_reg[1]0__1_n_108 ,\d_reg[1]0__1_n_109 ,\d_reg[1]0__1_n_110 ,\d_reg[1]0__1_n_111 ,\d_reg[1]0__1_n_112 ,\d_reg[1]0__1_n_113 ,\d_reg[1]0__1_n_114 ,\d_reg[1]0__1_n_115 ,\d_reg[1]0__1_n_116 ,\d_reg[1]0__1_n_117 ,\d_reg[1]0__1_n_118 ,\d_reg[1]0__1_n_119 ,\d_reg[1]0__1_n_120 ,\d_reg[1]0__1_n_121 ,\d_reg[1]0__1_n_122 ,\d_reg[1]0__1_n_123 ,\d_reg[1]0__1_n_124 ,\d_reg[1]0__1_n_125 ,\d_reg[1]0__1_n_126 ,\d_reg[1]0__1_n_127 ,\d_reg[1]0__1_n_128 ,\d_reg[1]0__1_n_129 ,\d_reg[1]0__1_n_130 ,\d_reg[1]0__1_n_131 ,\d_reg[1]0__1_n_132 ,\d_reg[1]0__1_n_133 ,\d_reg[1]0__1_n_134 ,\d_reg[1]0__1_n_135 ,\d_reg[1]0__1_n_136 ,\d_reg[1]0__1_n_137 ,\d_reg[1]0__1_n_138 ,\d_reg[1]0__1_n_139 ,\d_reg[1]0__1_n_140 ,\d_reg[1]0__1_n_141 ,\d_reg[1]0__1_n_142 ,\d_reg[1]0__1_n_143 ,\d_reg[1]0__1_n_144 ,\d_reg[1]0__1_n_145 ,\d_reg[1]0__1_n_146 ,\d_reg[1]0__1_n_147 ,\d_reg[1]0__1_n_148 ,\d_reg[1]0__1_n_149 ,\d_reg[1]0__1_n_150 ,\d_reg[1]0__1_n_151 ,\d_reg[1]0__1_n_152 ,\d_reg[1]0__1_n_153 }),
        .RSTA(RSTA),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(RSTA),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_1 
       (.I0(g0_b16_n_0),
        .I1(g1_b16_n_0),
        .O(\d_reg[1]0_i_1_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_10 
       (.I0(g0_b7_n_0),
        .I1(g1_b7_n_0),
        .O(\d_reg[1]0_i_10_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_10__0 
       (.I0(g0_b21_n_0),
        .I1(g1_b21_n_0),
        .O(\d_reg[1]0_i_10__0_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_11 
       (.I0(g0_b6_n_0),
        .I1(g1_b6_n_0),
        .O(\d_reg[1]0_i_11_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_11__0 
       (.I0(g0_b20_n_0),
        .I1(g1_b20_n_0),
        .O(\d_reg[1]0_i_11__0_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_12 
       (.I0(g0_b5_n_0),
        .I1(g1_b5_n_0),
        .O(\d_reg[1]0_i_12_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_12__0 
       (.I0(g0_b19_n_0),
        .I1(g1_b19_n_0),
        .O(\d_reg[1]0_i_12__0_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_13 
       (.I0(g0_b4_n_0),
        .I1(g1_b4_n_0),
        .O(\d_reg[1]0_i_13_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_13__0 
       (.I0(g0_b18_n_0),
        .I1(g1_b18_n_0),
        .O(\d_reg[1]0_i_13__0_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_14 
       (.I0(g0_b3_n_0),
        .I1(g1_b3_n_0),
        .O(\d_reg[1]0_i_14_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_14__0 
       (.I0(g0_b17_n_0),
        .I1(g1_b17_n_0),
        .O(\d_reg[1]0_i_14__0_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_15 
       (.I0(g0_b2_n_0),
        .I1(g1_b2_n_0),
        .O(\d_reg[1]0_i_15_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_16 
       (.I0(g0_b1_n_0),
        .I1(g1_b1_n_0),
        .O(\d_reg[1]0_i_16_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_17 
       (.I0(g0_b0_n_0),
        .I1(g1_b0_n_0),
        .O(\d_reg[1]0_i_17_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \d_reg[1]0_i_1__0 
       (.I0(g0_b30_n_0),
        .I1(ARG[29]),
        .O(\d_reg[1]0_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_2 
       (.I0(g0_b15_n_0),
        .I1(g1_b15_n_0),
        .O(\d_reg[1]0_i_2_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_2__0 
       (.I0(g0_b29_n_0),
        .I1(g1_b29_n_0),
        .O(\d_reg[1]0_i_2__0_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_3 
       (.I0(g0_b14_n_0),
        .I1(g1_b14_n_0),
        .O(\d_reg[1]0_i_3_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_3__0 
       (.I0(g0_b28_n_0),
        .I1(g1_b28_n_0),
        .O(\d_reg[1]0_i_3__0_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_4 
       (.I0(g0_b13_n_0),
        .I1(g1_b13_n_0),
        .O(\d_reg[1]0_i_4_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_4__0 
       (.I0(g0_b27_n_0),
        .I1(g1_b27_n_0),
        .O(\d_reg[1]0_i_4__0_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_5 
       (.I0(g0_b12_n_0),
        .I1(g1_b12_n_0),
        .O(\d_reg[1]0_i_5_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_5__0 
       (.I0(g0_b26_n_0),
        .I1(g1_b26_n_0),
        .O(\d_reg[1]0_i_5__0_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_6 
       (.I0(g0_b11_n_0),
        .I1(g1_b11_n_0),
        .O(\d_reg[1]0_i_6_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_6__0 
       (.I0(g0_b25_n_0),
        .I1(g1_b25_n_0),
        .O(\d_reg[1]0_i_6__0_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_7 
       (.I0(g0_b10_n_0),
        .I1(g1_b10_n_0),
        .O(\d_reg[1]0_i_7_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_7__0 
       (.I0(g0_b24_n_0),
        .I1(g1_b24_n_0),
        .O(\d_reg[1]0_i_7__0_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_8 
       (.I0(g0_b9_n_0),
        .I1(g1_b9_n_0),
        .O(\d_reg[1]0_i_8_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_8__0 
       (.I0(g0_b23_n_0),
        .I1(g1_b23_n_0),
        .O(\d_reg[1]0_i_8__0_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_9 
       (.I0(g0_b8_n_0),
        .I1(g1_b8_n_0),
        .O(\d_reg[1]0_i_9_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \d_reg[1]0_i_9__0 
       (.I0(g0_b22_n_0),
        .I1(g1_b22_n_0),
        .O(\d_reg[1]0_i_9__0_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDEB9084E8B6103E1)) 
    g0_b0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF6F69D2D1516A032)) 
    g0_b0__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b0__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h32DD4F9B81474F09)) 
    g0_b1
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h870AF8C93B8F9A51)) 
    g0_b10
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h56EB65F4A75C6A20)) 
    g0_b10__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b10__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h70B3DADD9F778EC1)) 
    g0_b11
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB76CEC98CA7A3B70)) 
    g0_b11__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b11__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0E58EEEF502E1CE5)) 
    g0_b12
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEAC9E58CE945F2D7)) 
    g0_b12__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b12__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF883FCAADDA4D1DD)) 
    g0_b13
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBAEC1E1E4BC27D19)) 
    g0_b13__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b13__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h516935F9082D45D5)) 
    g0_b14
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA15157A6EF9433B5)) 
    g0_b14__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b14__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAC58B5D88970603D)) 
    g0_b15
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b15_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB794CD3CCB2B2D73)) 
    g0_b15__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b15__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEDF4A812FFDB826D)) 
    g0_b16
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h767F0FA410779E5A)) 
    g0_b16__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b16__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2AEE4BE305DB325D)) 
    g0_b17
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b17_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE688872ADB6319FA)) 
    g0_b17__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b17__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF46C6B30CFAAD33D)) 
    g0_b18
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b18_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB9AFA88E666B5A27)) 
    g0_b18__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b18__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBD67C9E12DBD2A31)) 
    g0_b19
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b19_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h95306531D46666BE)) 
    g0_b19__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b19__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5AA4008B6CB91802)) 
    g0_b1__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0962CD28DDBC0AE1)) 
    g0_b2
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966288BF4CC5ED49)) 
    g0_b20
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8C9549C032CB8194)) 
    g0_b20__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b20__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h279E5D3F26FCB0D1)) 
    g0_b21
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD6D98E000E26AAD8)) 
    g0_b21__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b21__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3801C495B7039561)) 
    g0_b22
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE71E0FFFFE1E664A)) 
    g0_b22__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b22__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFFC38C92AAD981)) 
    g0_b23
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b23_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAD4AA55554AB4B6C)) 
    g0_b23__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b23__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h95556AD6DB331E01)) 
    g0_b24
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b24_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9CC663333266D925)) 
    g0_b24__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b24__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8CCCD9B249694AAB)) 
    g0_b25
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b25_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h83C1E0F0F1E1C71C)) 
    g0_b25__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b25__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7C3C3871C718C667)) 
    g0_b26
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b26_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7FC01FF00FE03F03)) 
    g0_b26__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b26__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFC03F80FC0F83E1F)) 
    g0_b27
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b27_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h003FFFF0001FFF00)) 
    g0_b27__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b27__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h03FFF8003FF801FF)) 
    g0_b28
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b28_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE03)) 
    g0_b28__0
       (.I0(ARG[25]),
        .I1(ARG[26]),
        .I2(ARG[27]),
        .I3(ARG[28]),
        .O(g0_b28__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF8000007FFFF)) 
    g0_b29
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b29_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h000001FF)) 
    g0_b29__0
       (.I0(ARG[25]),
        .I1(ARG[26]),
        .I2(ARG[27]),
        .I3(ARG[28]),
        .I4(ARG[29]),
        .O(g0_b29__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h66805AAD644AA059)) 
    g0_b2__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h394A3C90DBCD2B59)) 
    g0_b3
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000007FFFFFFFFFF)) 
    g0_b30
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b30_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9777E845E298C5A4)) 
    g0_b3__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h24ED2C5EB7370559)) 
    g0_b4
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h874AE5A699AAA4E9)) 
    g0_b4__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88F44BA7824BEC2D)) 
    g0_b5
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h91CB0D7B95C9D80B)) 
    g0_b5__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b5__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA3D86ED060390A9)) 
    g0_b6
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBB89793914129BF2)) 
    g0_b6__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b6__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h297A1098E599AD11)) 
    g0_b7
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h84CAEE993EAC8F24)) 
    g0_b7__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b7__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4035990796FC7E69)) 
    g0_b8
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3F0CCFBBA8C1AE83)) 
    g0_b8__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b8__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4AD2DC12E14CB3B1)) 
    g0_b9
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8B40BCAC278E3163)) 
    g0_b9__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g0_b9__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30A6DA0FFBC8AFF7)) 
    g1_b0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h604DF8B4C2E2050A)) 
    g1_b0__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b0__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5ED66BF04C2DE535)) 
    g1_b1
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h570A8F8473FE22AA)) 
    g1_b10
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h37D4C03AE05ABC44)) 
    g1_b10__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b10__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0C480B440E8C735D)) 
    g1_b11
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1CEC73AE8A03461D)) 
    g1_b11__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b11__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h247F5523CBD17FC6)) 
    g1_b12
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5D3A47CE15BC21BC)) 
    g1_b12__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b12__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h15E2C8257F4801BC)) 
    g1_b13
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h50773AA4F7198E83)) 
    g1_b13__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b13__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0E3AF6CCD1F6FF1B)) 
    g1_b14
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2450566258A5B94C)) 
    g1_b14__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b14__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h57ED893A53BA00A4)) 
    g1_b15
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b15_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h60A9FD2D060FF6E1)) 
    g1_b15__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b15__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h54D636DD8D7CAAC2)) 
    g1_b16
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3D1088A776EDB6C7)) 
    g1_b16__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b16__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1076E38D8D66AA98)) 
    g1_b17
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b17_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h160AFADD8CE6667D)) 
    g1_b17__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b17__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h382641065396220E)) 
    g1_b18
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b18_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0D5306560248137C)) 
    g1_b18__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b18__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0AB9D5FD60A67251)) 
    g1_b19
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b19_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0336AB67FE255B83)) 
    g1_b19__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b19__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2A3724FD8D844558)) 
    g1_b1__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h510765653CC63933)) 
    g1_b2
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h066A99FCD539E89F)) 
    g1_b20
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00F1992D54B663FF)) 
    g1_b20__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b20__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h01E64B5699C019B5)) 
    g1_b21
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000F871CCD92D6AA)) 
    g1_b21__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b21__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001E38CDB4AAAD26)) 
    g1_b22
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h55552A5696DB64CC)) 
    g1_b22__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b22__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5554AD6926CCCE38)) 
    g1_b23
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b23_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h333366CDB2492DA5)) 
    g1_b23__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b23__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h333264DB6DA5A56A)) 
    g1_b24
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b24_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0F0F1E3C71C71C63)) 
    g1_b24__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b24__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0F0E1C38E39C6319)) 
    g1_b25
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b25_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FF01FC0FC0FC1F)) 
    g1_b25__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b25__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FE03F81F83E0F8)) 
    g1_b26
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b26_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00FE07E0)) 
    g1_b26__0
       (.I0(ARG[24]),
        .I1(ARG[25]),
        .I2(ARG[26]),
        .I3(ARG[27]),
        .I4(ARG[28]),
        .O(g1_b26__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0001FFF8007FE007)) 
    g1_b27
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b27_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0001FFE0)) 
    g1_b27__0
       (.I0(ARG[24]),
        .I1(ARG[25]),
        .I2(ARG[26]),
        .I3(ARG[27]),
        .I4(ARG[28]),
        .O(g1_b27__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000007FFFFE000)) 
    g1_b28
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b28_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000001F)) 
    g1_b28__0
       (.I0(ARG[24]),
        .I1(ARG[25]),
        .I2(ARG[26]),
        .I3(ARG[27]),
        .I4(ARG[28]),
        .O(g1_b28__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000001FFF)) 
    g1_b29
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b29_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6EEEC6AFE0335345)) 
    g1_b2__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5839CD07B1AFF3A9)) 
    g1_b3
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5D9DD7108429BF19)) 
    g1_b3__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1F52631DF9CCA1CE)) 
    g1_b4
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h359B568D6B11E250)) 
    g1_b4__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1E735270AF024B74)) 
    g1_b5
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5379890C8ADB8455)) 
    g1_b5__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b5__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h25E257570113710A)) 
    g1_b6
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h65C4FB6C470B195F)) 
    g1_b6__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b6__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4D451478CE575CDC)) 
    g1_b7
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4AE8A388692F954A)) 
    g1_b7__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b7__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0D373BB1760DEDB7)) 
    g1_b8
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h402DD45480D4FF49)) 
    g1_b8__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b8__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h12325E760D35B9B9)) 
    g1_b9
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3861F94D8100D5AF)) 
    g1_b9__0
       (.I0(ARG[23]),
        .I1(ARG[24]),
        .I2(ARG[25]),
        .I3(ARG[26]),
        .I4(ARG[27]),
        .I5(ARG[28]),
        .O(g1_b9__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][0]_i_10 
       (.I0(\n_reg[3]0__2_n_97 ),
        .I1(\n_reg[3]0_n_97 ),
        .O(n));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][0]_i_11 
       (.I0(\n_reg[3]0__2_n_98 ),
        .I1(\n_reg[3]0_n_98 ),
        .O(\n[3][0]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][0]_i_13 
       (.I0(\n_reg[3]0__2_n_99 ),
        .I1(\n_reg[3]0_n_99 ),
        .O(\n[3][0]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][0]_i_14 
       (.I0(\n_reg[3]0__2_n_100 ),
        .I1(\n_reg[3]0_n_100 ),
        .O(\n[3][0]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][0]_i_15 
       (.I0(\n_reg[3]0__2_n_101 ),
        .I1(\n_reg[3]0_n_101 ),
        .O(\n[3][0]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][0]_i_16 
       (.I0(\n_reg[3]0__2_n_102 ),
        .I1(\n_reg[3]0_n_102 ),
        .O(\n[3][0]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][0]_i_17 
       (.I0(\n_reg[3]0__2_n_103 ),
        .I1(\n_reg[3]0_n_103 ),
        .O(\n[3][0]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][0]_i_18 
       (.I0(\n_reg[3]0__2_n_104 ),
        .I1(\n_reg[3]0_n_104 ),
        .O(\n[3][0]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][0]_i_19 
       (.I0(\n_reg[3]0__2_n_105 ),
        .I1(\n_reg[3]0_n_105 ),
        .O(\n[3][0]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][0]_i_3 
       (.I0(\n_reg[3]0__2_n_91 ),
        .I1(\n_reg[3]0_n_91 ),
        .O(\n[3][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][0]_i_4 
       (.I0(\n_reg[3]0__2_n_92 ),
        .I1(\n_reg[3]0_n_92 ),
        .O(\n[3][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][0]_i_5 
       (.I0(\n_reg[3]0__2_n_93 ),
        .I1(\n_reg[3]0_n_93 ),
        .O(\n[3][0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][0]_i_6 
       (.I0(\n_reg[3]0__2_n_94 ),
        .I1(\n_reg[3]0_n_94 ),
        .O(\n[3][0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][0]_i_8 
       (.I0(\n_reg[3]0__2_n_95 ),
        .I1(\n_reg[3]0_n_95 ),
        .O(\n[3][0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][0]_i_9 
       (.I0(\n_reg[3]0__2_n_96 ),
        .I1(\n_reg[3]0_n_96 ),
        .O(\n[3][0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][12]_i_2 
       (.I0(\n_reg[3]0__2_n_79 ),
        .I1(\n_reg[3]0__0_n_96 ),
        .O(\n[3][12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][12]_i_3 
       (.I0(\n_reg[3]0__2_n_80 ),
        .I1(\n_reg[3]0__0_n_97 ),
        .O(\n[3][12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][12]_i_4 
       (.I0(\n_reg[3]0__2_n_81 ),
        .I1(\n_reg[3]0__0_n_98 ),
        .O(\n[3][12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][12]_i_5 
       (.I0(\n_reg[3]0__2_n_82 ),
        .I1(\n_reg[3]0__0_n_99 ),
        .O(\n[3][12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][16]_i_2 
       (.I0(\n_reg[3]0__2_n_75 ),
        .I1(\n_reg[3]0__0_n_92 ),
        .O(\n[3][16]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][16]_i_3 
       (.I0(\n_reg[3]0__2_n_76 ),
        .I1(\n_reg[3]0__0_n_93 ),
        .O(\n[3][16]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][16]_i_4 
       (.I0(\n_reg[3]0__2_n_77 ),
        .I1(\n_reg[3]0__0_n_94 ),
        .O(\n[3][16]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][16]_i_5 
       (.I0(\n_reg[3]0__2_n_78 ),
        .I1(\n_reg[3]0__0_n_95 ),
        .O(\n[3][16]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][20]_i_2 
       (.I0(\n_reg[3]0__2_n_71 ),
        .I1(\n_reg[3]0__0_n_88 ),
        .O(\n[3][20]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][20]_i_3 
       (.I0(\n_reg[3]0__2_n_72 ),
        .I1(\n_reg[3]0__0_n_89 ),
        .O(\n[3][20]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][20]_i_4 
       (.I0(\n_reg[3]0__2_n_73 ),
        .I1(\n_reg[3]0__0_n_90 ),
        .O(\n[3][20]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][20]_i_5 
       (.I0(\n_reg[3]0__2_n_74 ),
        .I1(\n_reg[3]0__0_n_91 ),
        .O(\n[3][20]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][24]_i_2 
       (.I0(\n_reg[3]0__2_n_67 ),
        .I1(\n_reg[3]0__0_n_84 ),
        .O(\n[3][24]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][24]_i_3 
       (.I0(\n_reg[3]0__2_n_68 ),
        .I1(\n_reg[3]0__0_n_85 ),
        .O(\n[3][24]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][24]_i_4 
       (.I0(\n_reg[3]0__2_n_69 ),
        .I1(\n_reg[3]0__0_n_86 ),
        .O(\n[3][24]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][24]_i_5 
       (.I0(\n_reg[3]0__2_n_70 ),
        .I1(\n_reg[3]0__0_n_87 ),
        .O(\n[3][24]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][28]_i_2 
       (.I0(\n_reg[3]0__2_n_63 ),
        .I1(\n_reg[3]0__0_n_80 ),
        .O(\n[3][28]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][28]_i_3 
       (.I0(\n_reg[3]0__2_n_64 ),
        .I1(\n_reg[3]0__0_n_81 ),
        .O(\n[3][28]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][28]_i_4 
       (.I0(\n_reg[3]0__2_n_65 ),
        .I1(\n_reg[3]0__0_n_82 ),
        .O(\n[3][28]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][28]_i_5 
       (.I0(\n_reg[3]0__2_n_66 ),
        .I1(\n_reg[3]0__0_n_83 ),
        .O(\n[3][28]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n[3][31]_i_1 
       (.I0(res),
        .O(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][31]_i_3 
       (.I0(\n_reg[3]0__2_n_60 ),
        .I1(\n_reg[3]0__0_n_77 ),
        .O(\n[3][31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][31]_i_4 
       (.I0(\n_reg[3]0__2_n_61 ),
        .I1(\n_reg[3]0__0_n_78 ),
        .O(\n[3][31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][31]_i_5 
       (.I0(\n_reg[3]0__2_n_62 ),
        .I1(\n_reg[3]0__0_n_79 ),
        .O(\n[3][31]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][4]_i_2 
       (.I0(\n_reg[3]0__2_n_87 ),
        .I1(\n_reg[3]0__0_n_104 ),
        .O(\n[3][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][4]_i_3 
       (.I0(\n_reg[3]0__2_n_88 ),
        .I1(\n_reg[3]0__0_n_105 ),
        .O(\n[3][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][4]_i_4 
       (.I0(\n_reg[3]0__2_n_89 ),
        .I1(\n_reg[3]0_n_89 ),
        .O(\n[3][4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][4]_i_5 
       (.I0(\n_reg[3]0__2_n_90 ),
        .I1(\n_reg[3]0_n_90 ),
        .O(\n[3][4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][8]_i_2 
       (.I0(\n_reg[3]0__2_n_83 ),
        .I1(\n_reg[3]0__0_n_100 ),
        .O(\n[3][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][8]_i_3 
       (.I0(\n_reg[3]0__2_n_84 ),
        .I1(\n_reg[3]0__0_n_101 ),
        .O(\n[3][8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][8]_i_4 
       (.I0(\n_reg[3]0__2_n_85 ),
        .I1(\n_reg[3]0__0_n_102 ),
        .O(\n[3][8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n[3][8]_i_5 
       (.I0(\n_reg[3]0__2_n_86 ),
        .I1(\n_reg[3]0__0_n_103 ),
        .O(\n[3][8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-10 {cell *THIS*} {string 16x18 4}}" *) 
  DSP48E1 #(
    .ACASCREG(1),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(1),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(1),
    .BREG(1),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \n_reg[1]0 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\n_reg[1]0_i_1_n_0 ,\n_reg[1]0_i_2_n_0 ,\n_reg[1]0_i_3_n_0 ,\n_reg[1]0_i_4_n_0 ,\n_reg[1]0_i_5_n_0 ,\n_reg[1]0_i_6_n_0 ,\n_reg[1]0_i_7_n_0 ,\n_reg[1]0_i_8_n_0 ,\n_reg[1]0_i_9_n_0 ,\n_reg[1]0_i_10_n_0 ,\n_reg[1]0_i_11_n_0 ,\n_reg[1]0_i_12_n_0 ,\n_reg[1]0_i_13_n_0 ,\n_reg[1]0_i_14_n_0 ,\n_reg[1]0_i_15_n_0 ,\n_reg[1]0_i_16_n_0 ,\n_reg[1]0_i_17_n_0 }),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,ARG[31:17]}),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const1>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const1>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\n_reg[1]0_n_58 ,\n_reg[1]0_n_59 ,\n_reg[1]0_n_60 ,\n_reg[1]0_n_61 ,\n_reg[1]0_n_62 ,\n_reg[1]0_n_63 ,\n_reg[1]0_n_64 ,\n_reg[1]0_n_65 ,\n_reg[1]0_n_66 ,\n_reg[1]0_n_67 ,\n_reg[1]0_n_68 ,\n_reg[1]0_n_69 ,\n_reg[1]0_n_70 ,\n_reg[1]0_n_71 ,\n_reg[1]0_n_72 ,\n_reg[1]0_n_73 ,\n_reg[1]0_n_74 ,\n_reg[1]0_n_75 ,\n_reg[1]0_n_76 ,\n_reg[1]0_n_77 ,\n_reg[1]0_n_78 ,\n_reg[1]0_n_79 ,\n_reg[1]0_n_80 ,\n_reg[1]0_n_81 ,\n_reg[1]0_n_82 ,\n_reg[1]0_n_83 ,\n_reg[1]0_n_84 ,\n_reg[1]0_n_85 ,\n_reg[1]0_n_86 ,\n_reg[1]0_n_87 ,\n_reg[1]0_n_88 ,\n_reg[1]0_n_89 ,\n_reg[1]0_n_90 ,\n_reg[1]0_n_91 ,\n_reg[1]0_n_92 ,\n_reg[1]0_n_93 ,\n_reg[1]0_n_94 ,\n_reg[1]0_n_95 ,\n_reg[1]0_n_96 ,\n_reg[1]0_n_97 ,\n_reg[1]0_n_98 ,\n_reg[1]0_n_99 ,\n_reg[1]0_n_100 ,\n_reg[1]0_n_101 ,\n_reg[1]0_n_102 ,\n_reg[1]0_n_103 ,\n_reg[1]0_n_104 ,\n_reg[1]0_n_105 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .PCOUT({\n_reg[1]0_n_106 ,\n_reg[1]0_n_107 ,\n_reg[1]0_n_108 ,\n_reg[1]0_n_109 ,\n_reg[1]0_n_110 ,\n_reg[1]0_n_111 ,\n_reg[1]0_n_112 ,\n_reg[1]0_n_113 ,\n_reg[1]0_n_114 ,\n_reg[1]0_n_115 ,\n_reg[1]0_n_116 ,\n_reg[1]0_n_117 ,\n_reg[1]0_n_118 ,\n_reg[1]0_n_119 ,\n_reg[1]0_n_120 ,\n_reg[1]0_n_121 ,\n_reg[1]0_n_122 ,\n_reg[1]0_n_123 ,\n_reg[1]0_n_124 ,\n_reg[1]0_n_125 ,\n_reg[1]0_n_126 ,\n_reg[1]0_n_127 ,\n_reg[1]0_n_128 ,\n_reg[1]0_n_129 ,\n_reg[1]0_n_130 ,\n_reg[1]0_n_131 ,\n_reg[1]0_n_132 ,\n_reg[1]0_n_133 ,\n_reg[1]0_n_134 ,\n_reg[1]0_n_135 ,\n_reg[1]0_n_136 ,\n_reg[1]0_n_137 ,\n_reg[1]0_n_138 ,\n_reg[1]0_n_139 ,\n_reg[1]0_n_140 ,\n_reg[1]0_n_141 ,\n_reg[1]0_n_142 ,\n_reg[1]0_n_143 ,\n_reg[1]0_n_144 ,\n_reg[1]0_n_145 ,\n_reg[1]0_n_146 ,\n_reg[1]0_n_147 ,\n_reg[1]0_n_148 ,\n_reg[1]0_n_149 ,\n_reg[1]0_n_150 ,\n_reg[1]0_n_151 ,\n_reg[1]0_n_152 ,\n_reg[1]0_n_153 }),
        .RSTA(RSTA),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(RSTA),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-10 {cell *THIS*} {string 16x16 4}}" *) 
  DSP48E1 #(
    .ACASCREG(1),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(1),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(1),
    .BREG(1),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \n_reg[1]0__0 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,ARG[31:17]}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,g0_b29__0_n_0,\n_reg[1]0_i_1__0_n_0 ,\n_reg[1]0_i_2__0_n_0 ,\n_reg[1]0_i_3__0_n_0 ,\n_reg[1]0_i_4__0_n_0 ,\n_reg[1]0_i_5__0_n_0 ,\n_reg[1]0_i_6__0_n_0 ,\n_reg[1]0_i_7__0_n_0 ,\n_reg[1]0_i_8__0_n_0 ,\n_reg[1]0_i_9__0_n_0 ,\n_reg[1]0_i_10__0_n_0 ,\n_reg[1]0_i_11__0_n_0 ,\n_reg[1]0_i_12__0_n_0 }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const1>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const1>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P(n_reg),
        .PCIN({\n_reg[1]0_n_106 ,\n_reg[1]0_n_107 ,\n_reg[1]0_n_108 ,\n_reg[1]0_n_109 ,\n_reg[1]0_n_110 ,\n_reg[1]0_n_111 ,\n_reg[1]0_n_112 ,\n_reg[1]0_n_113 ,\n_reg[1]0_n_114 ,\n_reg[1]0_n_115 ,\n_reg[1]0_n_116 ,\n_reg[1]0_n_117 ,\n_reg[1]0_n_118 ,\n_reg[1]0_n_119 ,\n_reg[1]0_n_120 ,\n_reg[1]0_n_121 ,\n_reg[1]0_n_122 ,\n_reg[1]0_n_123 ,\n_reg[1]0_n_124 ,\n_reg[1]0_n_125 ,\n_reg[1]0_n_126 ,\n_reg[1]0_n_127 ,\n_reg[1]0_n_128 ,\n_reg[1]0_n_129 ,\n_reg[1]0_n_130 ,\n_reg[1]0_n_131 ,\n_reg[1]0_n_132 ,\n_reg[1]0_n_133 ,\n_reg[1]0_n_134 ,\n_reg[1]0_n_135 ,\n_reg[1]0_n_136 ,\n_reg[1]0_n_137 ,\n_reg[1]0_n_138 ,\n_reg[1]0_n_139 ,\n_reg[1]0_n_140 ,\n_reg[1]0_n_141 ,\n_reg[1]0_n_142 ,\n_reg[1]0_n_143 ,\n_reg[1]0_n_144 ,\n_reg[1]0_n_145 ,\n_reg[1]0_n_146 ,\n_reg[1]0_n_147 ,\n_reg[1]0_n_148 ,\n_reg[1]0_n_149 ,\n_reg[1]0_n_150 ,\n_reg[1]0_n_151 ,\n_reg[1]0_n_152 ,\n_reg[1]0_n_153 }),
        .RSTA(RSTA),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(RSTA),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-10 {cell *THIS*} {string 18x18 4}}" *) 
  DSP48E1 #(
    .ACASCREG(1),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(1),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(1),
    .BREG(1),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \n_reg[1]0__1 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,ARG[16:0]}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\n_reg[1]0_i_1_n_0 ,\n_reg[1]0_i_2_n_0 ,\n_reg[1]0_i_3_n_0 ,\n_reg[1]0_i_4_n_0 ,\n_reg[1]0_i_5_n_0 ,\n_reg[1]0_i_6_n_0 ,\n_reg[1]0_i_7_n_0 ,\n_reg[1]0_i_8_n_0 ,\n_reg[1]0_i_9_n_0 ,\n_reg[1]0_i_10_n_0 ,\n_reg[1]0_i_11_n_0 ,\n_reg[1]0_i_12_n_0 ,\n_reg[1]0_i_13_n_0 ,\n_reg[1]0_i_14_n_0 ,\n_reg[1]0_i_15_n_0 ,\n_reg[1]0_i_16_n_0 ,\n_reg[1]0_i_17_n_0 }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const1>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const1>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\n_reg[1]0__1_n_58 ,\n_reg[1]0__1_n_59 ,\n_reg[1]0__1_n_60 ,\n_reg[1]0__1_n_61 ,\n_reg[1]0__1_n_62 ,\n_reg[1]0__1_n_63 ,\n_reg[1]0__1_n_64 ,\n_reg[1]0__1_n_65 ,\n_reg[1]0__1_n_66 ,\n_reg[1]0__1_n_67 ,\n_reg[1]0__1_n_68 ,\n_reg[1]0__1_n_69 ,\n_reg[1]0__1_n_70 ,\n_reg[1]0__1_n_71 ,\n_reg[1]0__1_n_72 ,\n_reg[1]0__1_n_73 ,\n_reg[1]0__1_n_74 ,\n_reg[1]0__1_n_75 ,\n_reg[1]0__1_n_76 ,\n_reg[1]0__1_n_77 ,\n_reg[1]0__1_n_78 ,\n_reg[1]0__1_n_79 ,\n_reg[1]0__1_n_80 ,\n_reg[1]0__1_n_81 ,\n_reg[1]0__1_n_82 ,\n_reg[1]0__1_n_83 ,\n_reg[1]0__1_n_84 ,\n_reg[1]0__1_n_85 ,\n_reg[1]0__1_n_86 ,\n_reg[1]0__1_n_87 ,\n_reg[1]0__1_n_88 ,\n_reg[1]0__1_n_89 ,\n_reg[1]0__1_n_90 ,\n_reg[1]0__1_n_91 ,\n_reg[1]0__1_n_92 ,\n_reg[1]0__1_n_93 ,\n_reg[1]0__1_n_94 ,\n_reg[1]0__1_n_95 ,\n_reg[1]0__1_n_96 ,\n_reg[1]0__1_n_97 ,\n_reg[1]0__1_n_98 ,\n_reg[1]0__1_n_99 ,\n_reg[1]0__1_n_100 ,\n_reg[1]0__1_n_101 ,\n_reg[1]0__1_n_102 ,\n_reg[1]0__1_n_103 ,\n_reg[1]0__1_n_104 ,\n_reg[1]0__1_n_105 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .PCOUT({\n_reg[1]0__1_n_106 ,\n_reg[1]0__1_n_107 ,\n_reg[1]0__1_n_108 ,\n_reg[1]0__1_n_109 ,\n_reg[1]0__1_n_110 ,\n_reg[1]0__1_n_111 ,\n_reg[1]0__1_n_112 ,\n_reg[1]0__1_n_113 ,\n_reg[1]0__1_n_114 ,\n_reg[1]0__1_n_115 ,\n_reg[1]0__1_n_116 ,\n_reg[1]0__1_n_117 ,\n_reg[1]0__1_n_118 ,\n_reg[1]0__1_n_119 ,\n_reg[1]0__1_n_120 ,\n_reg[1]0__1_n_121 ,\n_reg[1]0__1_n_122 ,\n_reg[1]0__1_n_123 ,\n_reg[1]0__1_n_124 ,\n_reg[1]0__1_n_125 ,\n_reg[1]0__1_n_126 ,\n_reg[1]0__1_n_127 ,\n_reg[1]0__1_n_128 ,\n_reg[1]0__1_n_129 ,\n_reg[1]0__1_n_130 ,\n_reg[1]0__1_n_131 ,\n_reg[1]0__1_n_132 ,\n_reg[1]0__1_n_133 ,\n_reg[1]0__1_n_134 ,\n_reg[1]0__1_n_135 ,\n_reg[1]0__1_n_136 ,\n_reg[1]0__1_n_137 ,\n_reg[1]0__1_n_138 ,\n_reg[1]0__1_n_139 ,\n_reg[1]0__1_n_140 ,\n_reg[1]0__1_n_141 ,\n_reg[1]0__1_n_142 ,\n_reg[1]0__1_n_143 ,\n_reg[1]0__1_n_144 ,\n_reg[1]0__1_n_145 ,\n_reg[1]0__1_n_146 ,\n_reg[1]0__1_n_147 ,\n_reg[1]0__1_n_148 ,\n_reg[1]0__1_n_149 ,\n_reg[1]0__1_n_150 ,\n_reg[1]0__1_n_151 ,\n_reg[1]0__1_n_152 ,\n_reg[1]0__1_n_153 }),
        .RSTA(RSTA),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(RSTA),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-10 {cell *THIS*} {string 18x16 4}}" *) 
  DSP48E1 #(
    .ACASCREG(1),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(1),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(1),
    .BREG(1),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \n_reg[1]0__2 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,ARG[16:0]}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,g0_b29__0_n_0,\n_reg[1]0_i_1__0_n_0 ,\n_reg[1]0_i_2__0_n_0 ,\n_reg[1]0_i_3__0_n_0 ,\n_reg[1]0_i_4__0_n_0 ,\n_reg[1]0_i_5__0_n_0 ,\n_reg[1]0_i_6__0_n_0 ,\n_reg[1]0_i_7__0_n_0 ,\n_reg[1]0_i_8__0_n_0 ,\n_reg[1]0_i_9__0_n_0 ,\n_reg[1]0_i_10__0_n_0 ,\n_reg[1]0_i_11__0_n_0 ,\n_reg[1]0_i_12__0_n_0 }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const1>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const1>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\n_reg[1]0__2_n_58 ,\n_reg[1]0__2_n_59 ,\n_reg[1]0__2_n_60 ,\n_reg[1]0__2_n_61 ,\n_reg[1]0__2_n_62 ,\n_reg[1]0__2_n_63 ,\n_reg[1]0__2_n_64 ,\n_reg[1]0__2_n_65 ,\n_reg[1]0__2_n_66 ,\n_reg[1]0__2_n_67 ,\n_reg[1]0__2_n_68 ,\n_reg[1]0__2_n_69 ,\n_reg[1]0__2_n_70 ,\n_reg[1]0__2_n_71 ,\n_reg[1]0__2_n_72 ,\n_reg[1]0__2_n_73 ,\n_reg[1]0__2_n_74 ,\n_reg[1]0__2_n_75 ,\n_reg[1]0__2_n_76 ,\n_reg[1]0__2_n_77 ,\n_reg[1]0__2_n_78 ,\n_reg[1]0__2_n_79 ,\n_reg[1]0__2_n_80 ,\n_reg[1]0__2_n_81 ,\n_reg[1]0__2_n_82 ,\n_reg[1]0__2_n_83 ,\n_reg[1]0__2_n_84 ,\n_reg[1]0__2_n_85 ,\n_reg[1]0__2_n_86 ,\n_reg[1]0__2_n_87 ,\n_reg[1]0__2_n_88 ,\n_reg[1]0__2_n_89 ,\n_reg[1]0__2_n_90 ,\n_reg[1]0__2_n_91 ,\n_reg[1]0__2_n_92 ,\n_reg[1]0__2_n_93 ,\n_reg[1]0__2_n_94 ,\n_reg[1]0__2_n_95 ,\n_reg[1]0__2_n_96 ,\n_reg[1]0__2_n_97 ,\n_reg[1]0__2_n_98 ,\n_reg[1]0__2_n_99 ,\n_reg[1]0__2_n_100 ,\n_reg[1]0__2_n_101 ,\n_reg[1]0__2_n_102 ,\n_reg[1]0__2_n_103 ,\n_reg[1]0__2_n_104 ,\n_reg[1]0__2_n_105 }),
        .PCIN({\n_reg[1]0__1_n_106 ,\n_reg[1]0__1_n_107 ,\n_reg[1]0__1_n_108 ,\n_reg[1]0__1_n_109 ,\n_reg[1]0__1_n_110 ,\n_reg[1]0__1_n_111 ,\n_reg[1]0__1_n_112 ,\n_reg[1]0__1_n_113 ,\n_reg[1]0__1_n_114 ,\n_reg[1]0__1_n_115 ,\n_reg[1]0__1_n_116 ,\n_reg[1]0__1_n_117 ,\n_reg[1]0__1_n_118 ,\n_reg[1]0__1_n_119 ,\n_reg[1]0__1_n_120 ,\n_reg[1]0__1_n_121 ,\n_reg[1]0__1_n_122 ,\n_reg[1]0__1_n_123 ,\n_reg[1]0__1_n_124 ,\n_reg[1]0__1_n_125 ,\n_reg[1]0__1_n_126 ,\n_reg[1]0__1_n_127 ,\n_reg[1]0__1_n_128 ,\n_reg[1]0__1_n_129 ,\n_reg[1]0__1_n_130 ,\n_reg[1]0__1_n_131 ,\n_reg[1]0__1_n_132 ,\n_reg[1]0__1_n_133 ,\n_reg[1]0__1_n_134 ,\n_reg[1]0__1_n_135 ,\n_reg[1]0__1_n_136 ,\n_reg[1]0__1_n_137 ,\n_reg[1]0__1_n_138 ,\n_reg[1]0__1_n_139 ,\n_reg[1]0__1_n_140 ,\n_reg[1]0__1_n_141 ,\n_reg[1]0__1_n_142 ,\n_reg[1]0__1_n_143 ,\n_reg[1]0__1_n_144 ,\n_reg[1]0__1_n_145 ,\n_reg[1]0__1_n_146 ,\n_reg[1]0__1_n_147 ,\n_reg[1]0__1_n_148 ,\n_reg[1]0__1_n_149 ,\n_reg[1]0__1_n_150 ,\n_reg[1]0__1_n_151 ,\n_reg[1]0__1_n_152 ,\n_reg[1]0__1_n_153 }),
        .RSTA(RSTA),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(RSTA),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_1 
       (.I0(g0_b16__0_n_0),
        .I1(g1_b16__0_n_0),
        .O(\n_reg[1]0_i_1_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_10 
       (.I0(g0_b7__0_n_0),
        .I1(g1_b7__0_n_0),
        .O(\n_reg[1]0_i_10_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_10__0 
       (.I0(g0_b19__0_n_0),
        .I1(g1_b19__0_n_0),
        .O(\n_reg[1]0_i_10__0_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_11 
       (.I0(g0_b6__0_n_0),
        .I1(g1_b6__0_n_0),
        .O(\n_reg[1]0_i_11_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_11__0 
       (.I0(g0_b18__0_n_0),
        .I1(g1_b18__0_n_0),
        .O(\n_reg[1]0_i_11__0_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_12 
       (.I0(g0_b5__0_n_0),
        .I1(g1_b5__0_n_0),
        .O(\n_reg[1]0_i_12_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_12__0 
       (.I0(g0_b17__0_n_0),
        .I1(g1_b17__0_n_0),
        .O(\n_reg[1]0_i_12__0_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_13 
       (.I0(g0_b4__0_n_0),
        .I1(g1_b4__0_n_0),
        .O(\n_reg[1]0_i_13_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_14 
       (.I0(g0_b3__0_n_0),
        .I1(g1_b3__0_n_0),
        .O(\n_reg[1]0_i_14_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_15 
       (.I0(g0_b2__0_n_0),
        .I1(g1_b2__0_n_0),
        .O(\n_reg[1]0_i_15_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_16 
       (.I0(g0_b1__0_n_0),
        .I1(g1_b1__0_n_0),
        .O(\n_reg[1]0_i_16_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_17 
       (.I0(g0_b0__0_n_0),
        .I1(g1_b0__0_n_0),
        .O(\n_reg[1]0_i_17_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \n_reg[1]0_i_1__0 
       (.I0(g0_b28__0_n_0),
        .I1(g1_b28__0_n_0),
        .I2(ARG[29]),
        .O(\n_reg[1]0_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_2 
       (.I0(g0_b15__0_n_0),
        .I1(g1_b15__0_n_0),
        .O(\n_reg[1]0_i_2_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_2__0 
       (.I0(g0_b27__0_n_0),
        .I1(g1_b27__0_n_0),
        .O(\n_reg[1]0_i_2__0_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_3 
       (.I0(g0_b14__0_n_0),
        .I1(g1_b14__0_n_0),
        .O(\n_reg[1]0_i_3_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_3__0 
       (.I0(g0_b26__0_n_0),
        .I1(g1_b26__0_n_0),
        .O(\n_reg[1]0_i_3__0_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_4 
       (.I0(g0_b13__0_n_0),
        .I1(g1_b13__0_n_0),
        .O(\n_reg[1]0_i_4_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_4__0 
       (.I0(g0_b25__0_n_0),
        .I1(g1_b25__0_n_0),
        .O(\n_reg[1]0_i_4__0_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_5 
       (.I0(g0_b12__0_n_0),
        .I1(g1_b12__0_n_0),
        .O(\n_reg[1]0_i_5_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_5__0 
       (.I0(g0_b24__0_n_0),
        .I1(g1_b24__0_n_0),
        .O(\n_reg[1]0_i_5__0_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_6 
       (.I0(g0_b11__0_n_0),
        .I1(g1_b11__0_n_0),
        .O(\n_reg[1]0_i_6_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_6__0 
       (.I0(g0_b23__0_n_0),
        .I1(g1_b23__0_n_0),
        .O(\n_reg[1]0_i_6__0_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_7 
       (.I0(g0_b10__0_n_0),
        .I1(g1_b10__0_n_0),
        .O(\n_reg[1]0_i_7_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_7__0 
       (.I0(g0_b22__0_n_0),
        .I1(g1_b22__0_n_0),
        .O(\n_reg[1]0_i_7__0_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_8 
       (.I0(g0_b9__0_n_0),
        .I1(g1_b9__0_n_0),
        .O(\n_reg[1]0_i_8_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_8__0 
       (.I0(g0_b21__0_n_0),
        .I1(g1_b21__0_n_0),
        .O(\n_reg[1]0_i_8__0_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_9 
       (.I0(g0_b8__0_n_0),
        .I1(g1_b8__0_n_0),
        .O(\n_reg[1]0_i_9_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \n_reg[1]0_i_9__0 
       (.I0(g0_b20__0_n_0),
        .I1(g1_b20__0_n_0),
        .O(\n_reg[1]0_i_9__0_n_0 ),
        .S(ARG[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-10 {cell *THIS*} {string 16x18 4}}" *) 
  DSP48E1 #(
    .ACASCREG(1),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(1),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(1),
    .BREG(1),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \n_reg[2]0 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\r_reg[1]0 [16:1],\d_next[1] [1]}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\n_next[1] [31:17]}),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const1>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const1>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\n_reg[2]0_n_58 ,\n_reg[2]0_n_59 ,\n_reg[2]0_n_60 ,\n_reg[2]0_n_61 ,\n_reg[2]0_n_62 ,\n_reg[2]0_n_63 ,\n_reg[2]0_n_64 ,\n_reg[2]0_n_65 ,\n_reg[2]0_n_66 ,\n_reg[2]0_n_67 ,\n_reg[2]0_n_68 ,\n_reg[2]0_n_69 ,\n_reg[2]0_n_70 ,\n_reg[2]0_n_71 ,\n_reg[2]0_n_72 ,\n_reg[2]0_n_73 ,\n_reg[2]0_n_74 ,\n_reg[2]0_n_75 ,\n_reg[2]0_n_76 ,\n_reg[2]0_n_77 ,\n_reg[2]0_n_78 ,\n_reg[2]0_n_79 ,\n_reg[2]0_n_80 ,\n_reg[2]0_n_81 ,\n_reg[2]0_n_82 ,\n_reg[2]0_n_83 ,\n_reg[2]0_n_84 ,\n_reg[2]0_n_85 ,\n_reg[2]0_n_86 ,\n_reg[2]0_n_87 ,\n_reg[2]0_n_88 ,\n_reg[2]0_n_89 ,\n_reg[2]0_n_90 ,\n_reg[2]0_n_91 ,\n_reg[2]0_n_92 ,\n_reg[2]0_n_93 ,\n_reg[2]0_n_94 ,\n_reg[2]0_n_95 ,\n_reg[2]0_n_96 ,\n_reg[2]0_n_97 ,\n_reg[2]0_n_98 ,\n_reg[2]0_n_99 ,\n_reg[2]0_n_100 ,\n_reg[2]0_n_101 ,\n_reg[2]0_n_102 ,\n_reg[2]0_n_103 ,\n_reg[2]0_n_104 ,\n_reg[2]0_n_105 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .PCOUT({\n_reg[2]0_n_106 ,\n_reg[2]0_n_107 ,\n_reg[2]0_n_108 ,\n_reg[2]0_n_109 ,\n_reg[2]0_n_110 ,\n_reg[2]0_n_111 ,\n_reg[2]0_n_112 ,\n_reg[2]0_n_113 ,\n_reg[2]0_n_114 ,\n_reg[2]0_n_115 ,\n_reg[2]0_n_116 ,\n_reg[2]0_n_117 ,\n_reg[2]0_n_118 ,\n_reg[2]0_n_119 ,\n_reg[2]0_n_120 ,\n_reg[2]0_n_121 ,\n_reg[2]0_n_122 ,\n_reg[2]0_n_123 ,\n_reg[2]0_n_124 ,\n_reg[2]0_n_125 ,\n_reg[2]0_n_126 ,\n_reg[2]0_n_127 ,\n_reg[2]0_n_128 ,\n_reg[2]0_n_129 ,\n_reg[2]0_n_130 ,\n_reg[2]0_n_131 ,\n_reg[2]0_n_132 ,\n_reg[2]0_n_133 ,\n_reg[2]0_n_134 ,\n_reg[2]0_n_135 ,\n_reg[2]0_n_136 ,\n_reg[2]0_n_137 ,\n_reg[2]0_n_138 ,\n_reg[2]0_n_139 ,\n_reg[2]0_n_140 ,\n_reg[2]0_n_141 ,\n_reg[2]0_n_142 ,\n_reg[2]0_n_143 ,\n_reg[2]0_n_144 ,\n_reg[2]0_n_145 ,\n_reg[2]0_n_146 ,\n_reg[2]0_n_147 ,\n_reg[2]0_n_148 ,\n_reg[2]0_n_149 ,\n_reg[2]0_n_150 ,\n_reg[2]0_n_151 ,\n_reg[2]0_n_152 ,\n_reg[2]0_n_153 }),
        .RSTA(RSTA),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(RSTA),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-10 {cell *THIS*} {string 16x16 4}}" *) 
  DSP48E1 #(
    .ACASCREG(1),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(1),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(1),
    .BREG(1),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \n_reg[2]0__0 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\n_next[1] [31:17]}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\r_reg[1]0 [31:17]}),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const1>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const1>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\n_reg[2]0__0_n_58 ,\n_reg[2]0__0_n_59 ,\n_reg[2]0__0_n_60 ,\n_reg[2]0__0_n_61 ,\n_reg[2]0__0_n_62 ,\n_reg[2]0__0_n_63 ,\n_reg[2]0__0_n_64 ,\n_reg[2]0__0_n_65 ,\n_reg[2]0__0_n_66 ,\n_reg[2]0__0_n_67 ,\n_reg[2]0__0_n_68 ,\n_reg[2]0__0_n_69 ,\n_reg[2]0__0_n_70 ,\n_reg[2]0__0_n_71 ,\n_reg[2]0__0_n_72 ,\n_reg[2]0__0_n_73 ,\n_reg[2]0__0_n_74 ,\n_reg[2]0__0_n_75 ,\n_reg[2]0__0_n_76 ,\n_reg[2]0__0_n_77 ,\n_reg[2]0__0_n_78 ,\n_reg[2]0__0_n_79 ,\n_reg[2]0__0_n_80 ,\n_reg[2]0__0_n_81 ,\n_reg[2]0__0_n_82 ,\n_reg[2]0__0_n_83 ,\n_reg[2]0__0_n_84 ,\n_reg[2]0__0_n_85 ,\n_reg[2]0__0_n_86 ,\n_reg[2]0__0_n_87 ,\n_reg[2]0__0_n_88 ,\n_reg[2]0__0_n_89 ,\n_reg[2]0__0_n_90 ,\n_reg[2]0__0_n_91 ,\n_reg[2]0__0_n_92 ,\n_reg[2]0__0_n_93 ,\n_reg[2]0__0_n_94 ,\n_reg[2]0__0_n_95 ,\n_reg[2]0__0_n_96 ,\n_reg[2]0__0_n_97 ,\n_reg[2]0__0_n_98 ,\n_reg[2]0__0_n_99 ,\n_reg[2]0__0_n_100 ,\n_reg[2]0__0_n_101 ,\n_reg[2]0__0_n_102 ,\n_reg[2]0__0_n_103 ,\n_reg[2]0__0_n_104 ,\n_reg[2]0__0_n_105 }),
        .PCIN({\n_reg[2]0_n_106 ,\n_reg[2]0_n_107 ,\n_reg[2]0_n_108 ,\n_reg[2]0_n_109 ,\n_reg[2]0_n_110 ,\n_reg[2]0_n_111 ,\n_reg[2]0_n_112 ,\n_reg[2]0_n_113 ,\n_reg[2]0_n_114 ,\n_reg[2]0_n_115 ,\n_reg[2]0_n_116 ,\n_reg[2]0_n_117 ,\n_reg[2]0_n_118 ,\n_reg[2]0_n_119 ,\n_reg[2]0_n_120 ,\n_reg[2]0_n_121 ,\n_reg[2]0_n_122 ,\n_reg[2]0_n_123 ,\n_reg[2]0_n_124 ,\n_reg[2]0_n_125 ,\n_reg[2]0_n_126 ,\n_reg[2]0_n_127 ,\n_reg[2]0_n_128 ,\n_reg[2]0_n_129 ,\n_reg[2]0_n_130 ,\n_reg[2]0_n_131 ,\n_reg[2]0_n_132 ,\n_reg[2]0_n_133 ,\n_reg[2]0_n_134 ,\n_reg[2]0_n_135 ,\n_reg[2]0_n_136 ,\n_reg[2]0_n_137 ,\n_reg[2]0_n_138 ,\n_reg[2]0_n_139 ,\n_reg[2]0_n_140 ,\n_reg[2]0_n_141 ,\n_reg[2]0_n_142 ,\n_reg[2]0_n_143 ,\n_reg[2]0_n_144 ,\n_reg[2]0_n_145 ,\n_reg[2]0_n_146 ,\n_reg[2]0_n_147 ,\n_reg[2]0_n_148 ,\n_reg[2]0_n_149 ,\n_reg[2]0_n_150 ,\n_reg[2]0_n_151 ,\n_reg[2]0_n_152 ,\n_reg[2]0_n_153 }),
        .RSTA(RSTA),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(RSTA),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-10 {cell *THIS*} {string 18x18 4}}" *) 
  DSP48E1 #(
    .ACASCREG(1),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(1),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(1),
    .BREG(1),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \n_reg[2]0__1 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\n_next[1] [16:0]}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ACOUT({\n_reg[2]0__1_n_24 ,\n_reg[2]0__1_n_25 ,\n_reg[2]0__1_n_26 ,\n_reg[2]0__1_n_27 ,\n_reg[2]0__1_n_28 ,\n_reg[2]0__1_n_29 ,\n_reg[2]0__1_n_30 ,\n_reg[2]0__1_n_31 ,\n_reg[2]0__1_n_32 ,\n_reg[2]0__1_n_33 ,\n_reg[2]0__1_n_34 ,\n_reg[2]0__1_n_35 ,\n_reg[2]0__1_n_36 ,\n_reg[2]0__1_n_37 ,\n_reg[2]0__1_n_38 ,\n_reg[2]0__1_n_39 ,\n_reg[2]0__1_n_40 ,\n_reg[2]0__1_n_41 ,\n_reg[2]0__1_n_42 ,\n_reg[2]0__1_n_43 ,\n_reg[2]0__1_n_44 ,\n_reg[2]0__1_n_45 ,\n_reg[2]0__1_n_46 ,\n_reg[2]0__1_n_47 ,\n_reg[2]0__1_n_48 ,\n_reg[2]0__1_n_49 ,\n_reg[2]0__1_n_50 ,\n_reg[2]0__1_n_51 ,\n_reg[2]0__1_n_52 ,\n_reg[2]0__1_n_53 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\r_reg[1]0 [16:1],\d_next[1] [1]}),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const1>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const1>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\n_reg[2]0__1_n_58 ,\n_reg[2]0__1_n_59 ,\n_reg[2]0__1_n_60 ,\n_reg[2]0__1_n_61 ,\n_reg[2]0__1_n_62 ,\n_reg[2]0__1_n_63 ,\n_reg[2]0__1_n_64 ,\n_reg[2]0__1_n_65 ,\n_reg[2]0__1_n_66 ,\n_reg[2]0__1_n_67 ,\n_reg[2]0__1_n_68 ,\n_reg[2]0__1_n_69 ,\n_reg[2]0__1_n_70 ,\n_reg[2]0__1_n_71 ,\n_reg[2]0__1_n_72 ,\n_reg[2]0__1_n_73 ,\n_reg[2]0__1_n_74 ,\n_reg[2]0__1_n_75 ,\n_reg[2]0__1_n_76 ,\n_reg[2]0__1_n_77 ,\n_reg[2]0__1_n_78 ,\n_reg[2]0__1_n_79 ,\n_reg[2]0__1_n_80 ,\n_reg[2]0__1_n_81 ,\n_reg[2]0__1_n_82 ,\n_reg[2]0__1_n_83 ,\n_reg[2]0__1_n_84 ,\n_reg[2]0__1_n_85 ,\n_reg[2]0__1_n_86 ,\n_reg[2]0__1_n_87 ,\n_reg[2]0__1_n_88 ,\n_reg[2]0__1_n_89 ,\n_reg[2]0__1_n_90 ,\n_reg[2]0__1_n_91 ,\n_reg[2]0__1_n_92 ,\n_reg[2]0__1_n_93 ,\n_reg[2]0__1_n_94 ,\n_reg[2]0__1_n_95 ,\n_reg[2]0__1_n_96 ,\n_reg[2]0__1_n_97 ,\n_reg[2]0__1_n_98 ,\n_reg[2]0__1_n_99 ,\n_reg[2]0__1_n_100 ,\n_reg[2]0__1_n_101 ,\n_reg[2]0__1_n_102 ,\n_reg[2]0__1_n_103 ,\n_reg[2]0__1_n_104 ,\n_reg[2]0__1_n_105 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .PCOUT({\n_reg[2]0__1_n_106 ,\n_reg[2]0__1_n_107 ,\n_reg[2]0__1_n_108 ,\n_reg[2]0__1_n_109 ,\n_reg[2]0__1_n_110 ,\n_reg[2]0__1_n_111 ,\n_reg[2]0__1_n_112 ,\n_reg[2]0__1_n_113 ,\n_reg[2]0__1_n_114 ,\n_reg[2]0__1_n_115 ,\n_reg[2]0__1_n_116 ,\n_reg[2]0__1_n_117 ,\n_reg[2]0__1_n_118 ,\n_reg[2]0__1_n_119 ,\n_reg[2]0__1_n_120 ,\n_reg[2]0__1_n_121 ,\n_reg[2]0__1_n_122 ,\n_reg[2]0__1_n_123 ,\n_reg[2]0__1_n_124 ,\n_reg[2]0__1_n_125 ,\n_reg[2]0__1_n_126 ,\n_reg[2]0__1_n_127 ,\n_reg[2]0__1_n_128 ,\n_reg[2]0__1_n_129 ,\n_reg[2]0__1_n_130 ,\n_reg[2]0__1_n_131 ,\n_reg[2]0__1_n_132 ,\n_reg[2]0__1_n_133 ,\n_reg[2]0__1_n_134 ,\n_reg[2]0__1_n_135 ,\n_reg[2]0__1_n_136 ,\n_reg[2]0__1_n_137 ,\n_reg[2]0__1_n_138 ,\n_reg[2]0__1_n_139 ,\n_reg[2]0__1_n_140 ,\n_reg[2]0__1_n_141 ,\n_reg[2]0__1_n_142 ,\n_reg[2]0__1_n_143 ,\n_reg[2]0__1_n_144 ,\n_reg[2]0__1_n_145 ,\n_reg[2]0__1_n_146 ,\n_reg[2]0__1_n_147 ,\n_reg[2]0__1_n_148 ,\n_reg[2]0__1_n_149 ,\n_reg[2]0__1_n_150 ,\n_reg[2]0__1_n_151 ,\n_reg[2]0__1_n_152 ,\n_reg[2]0__1_n_153 }),
        .RSTA(RSTA),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(RSTA),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-10 {cell *THIS*} {string 18x16 4}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("CASCADE"),
    .BCASCREG(1),
    .BREG(1),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \n_reg[2]0__2 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ACIN({\n_reg[2]0__1_n_24 ,\n_reg[2]0__1_n_25 ,\n_reg[2]0__1_n_26 ,\n_reg[2]0__1_n_27 ,\n_reg[2]0__1_n_28 ,\n_reg[2]0__1_n_29 ,\n_reg[2]0__1_n_30 ,\n_reg[2]0__1_n_31 ,\n_reg[2]0__1_n_32 ,\n_reg[2]0__1_n_33 ,\n_reg[2]0__1_n_34 ,\n_reg[2]0__1_n_35 ,\n_reg[2]0__1_n_36 ,\n_reg[2]0__1_n_37 ,\n_reg[2]0__1_n_38 ,\n_reg[2]0__1_n_39 ,\n_reg[2]0__1_n_40 ,\n_reg[2]0__1_n_41 ,\n_reg[2]0__1_n_42 ,\n_reg[2]0__1_n_43 ,\n_reg[2]0__1_n_44 ,\n_reg[2]0__1_n_45 ,\n_reg[2]0__1_n_46 ,\n_reg[2]0__1_n_47 ,\n_reg[2]0__1_n_48 ,\n_reg[2]0__1_n_49 ,\n_reg[2]0__1_n_50 ,\n_reg[2]0__1_n_51 ,\n_reg[2]0__1_n_52 ,\n_reg[2]0__1_n_53 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\r_reg[1]0 [31:17]}),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const1>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\n_reg[2]0__2_n_58 ,\n_reg[2]0__2_n_59 ,\n_reg[2]0__2_n_60 ,\n_reg[2]0__2_n_61 ,\n_reg[2]0__2_n_62 ,\n_reg[2]0__2_n_63 ,\n_reg[2]0__2_n_64 ,\n_reg[2]0__2_n_65 ,\n_reg[2]0__2_n_66 ,\n_reg[2]0__2_n_67 ,\n_reg[2]0__2_n_68 ,\n_reg[2]0__2_n_69 ,\n_reg[2]0__2_n_70 ,\n_reg[2]0__2_n_71 ,\n_reg[2]0__2_n_72 ,\n_reg[2]0__2_n_73 ,\n_reg[2]0__2_n_74 ,\n_reg[2]0__2_n_75 ,\n_reg[2]0__2_n_76 ,\n_reg[2]0__2_n_77 ,\n_reg[2]0__2_n_78 ,\n_reg[2]0__2_n_79 ,\n_reg[2]0__2_n_80 ,\n_reg[2]0__2_n_81 ,\n_reg[2]0__2_n_82 ,\n_reg[2]0__2_n_83 ,\n_reg[2]0__2_n_84 ,\n_reg[2]0__2_n_85 ,\n_reg[2]0__2_n_86 ,\n_reg[2]0__2_n_87 ,\n_reg[2]0__2_n_88 ,\n_reg[2]0__2_n_89 ,\n_reg[2]0__2_n_90 ,\n_reg[2]0__2_n_91 ,\n_reg[2]0__2_n_92 ,\n_reg[2]0__2_n_93 ,\n_reg[2]0__2_n_94 ,\n_reg[2]0__2_n_95 ,\n_reg[2]0__2_n_96 ,\n_reg[2]0__2_n_97 ,\n_reg[2]0__2_n_98 ,\n_reg[2]0__2_n_99 ,\n_reg[2]0__2_n_100 ,\n_reg[2]0__2_n_101 ,\n_reg[2]0__2_n_102 ,\n_reg[2]0__2_n_103 ,\n_reg[2]0__2_n_104 ,\n_reg[2]0__2_n_105 }),
        .PCIN({\n_reg[2]0__1_n_106 ,\n_reg[2]0__1_n_107 ,\n_reg[2]0__1_n_108 ,\n_reg[2]0__1_n_109 ,\n_reg[2]0__1_n_110 ,\n_reg[2]0__1_n_111 ,\n_reg[2]0__1_n_112 ,\n_reg[2]0__1_n_113 ,\n_reg[2]0__1_n_114 ,\n_reg[2]0__1_n_115 ,\n_reg[2]0__1_n_116 ,\n_reg[2]0__1_n_117 ,\n_reg[2]0__1_n_118 ,\n_reg[2]0__1_n_119 ,\n_reg[2]0__1_n_120 ,\n_reg[2]0__1_n_121 ,\n_reg[2]0__1_n_122 ,\n_reg[2]0__1_n_123 ,\n_reg[2]0__1_n_124 ,\n_reg[2]0__1_n_125 ,\n_reg[2]0__1_n_126 ,\n_reg[2]0__1_n_127 ,\n_reg[2]0__1_n_128 ,\n_reg[2]0__1_n_129 ,\n_reg[2]0__1_n_130 ,\n_reg[2]0__1_n_131 ,\n_reg[2]0__1_n_132 ,\n_reg[2]0__1_n_133 ,\n_reg[2]0__1_n_134 ,\n_reg[2]0__1_n_135 ,\n_reg[2]0__1_n_136 ,\n_reg[2]0__1_n_137 ,\n_reg[2]0__1_n_138 ,\n_reg[2]0__1_n_139 ,\n_reg[2]0__1_n_140 ,\n_reg[2]0__1_n_141 ,\n_reg[2]0__1_n_142 ,\n_reg[2]0__1_n_143 ,\n_reg[2]0__1_n_144 ,\n_reg[2]0__1_n_145 ,\n_reg[2]0__1_n_146 ,\n_reg[2]0__1_n_147 ,\n_reg[2]0__1_n_148 ,\n_reg[2]0__1_n_149 ,\n_reg[2]0__1_n_150 ,\n_reg[2]0__1_n_151 ,\n_reg[2]0__1_n_152 ,\n_reg[2]0__1_n_153 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(RSTA),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[2]0_i_1 
       (.CI(\n_reg[2]0_i_2_n_0 ),
        .CO({\n_reg[2]0_i_1_n_0 ,\n_reg[2]0_i_1_n_1 ,\n_reg[2]0_i_1_n_2 ,\n_reg[2]0_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[1]0__2_n_75 ,\n_reg[1]0__2_n_76 ,\n_reg[1]0__2_n_77 ,\n_reg[1]0__2_n_78 }),
        .O(\n_next[1] [16:13]),
        .S({\n_reg[2]0_i_6_n_0 ,\n_reg[2]0_i_7_n_0 ,\n_reg[2]0_i_8_n_0 ,\n_reg[2]0_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_10 
       (.I0(\n_reg[1]0__2_n_79 ),
        .I1(n_reg[9]),
        .O(\n_reg[2]0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_10__0 
       (.I0(\n_reg[1]0__2_n_65 ),
        .I1(n_reg[23]),
        .O(\n_reg[2]0_i_10__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_11 
       (.I0(\n_reg[1]0__2_n_80 ),
        .I1(n_reg[8]),
        .O(\n_reg[2]0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_11__0 
       (.I0(\n_reg[1]0__2_n_66 ),
        .I1(n_reg[22]),
        .O(\n_reg[2]0_i_11__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_12 
       (.I0(\n_reg[1]0__2_n_81 ),
        .I1(n_reg[7]),
        .O(\n_reg[2]0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_12__0 
       (.I0(\n_reg[1]0__2_n_67 ),
        .I1(n_reg[21]),
        .O(\n_reg[2]0_i_12__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_13 
       (.I0(\n_reg[1]0__2_n_82 ),
        .I1(n_reg[6]),
        .O(\n_reg[2]0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_13__0 
       (.I0(\n_reg[1]0__2_n_68 ),
        .I1(n_reg[20]),
        .O(\n_reg[2]0_i_13__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_14 
       (.I0(\n_reg[1]0__2_n_83 ),
        .I1(n_reg[5]),
        .O(\n_reg[2]0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_14__0 
       (.I0(\n_reg[1]0__2_n_69 ),
        .I1(n_reg[19]),
        .O(\n_reg[2]0_i_14__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_15 
       (.I0(\n_reg[1]0__2_n_84 ),
        .I1(n_reg[4]),
        .O(\n_reg[2]0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_15__0 
       (.I0(\n_reg[1]0__2_n_70 ),
        .I1(n_reg[18]),
        .O(\n_reg[2]0_i_15__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_16 
       (.I0(\n_reg[1]0__2_n_85 ),
        .I1(n_reg[3]),
        .O(\n_reg[2]0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_16__0 
       (.I0(\n_reg[1]0__2_n_71 ),
        .I1(n_reg[17]),
        .O(\n_reg[2]0_i_16__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_17 
       (.I0(\n_reg[1]0__2_n_86 ),
        .I1(n_reg[2]),
        .O(\n_reg[2]0_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_17__0 
       (.I0(\n_reg[1]0__2_n_72 ),
        .I1(n_reg[16]),
        .O(\n_reg[2]0_i_17__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_18 
       (.I0(\n_reg[1]0__2_n_87 ),
        .I1(n_reg[1]),
        .O(\n_reg[2]0_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_18__0 
       (.I0(\n_reg[1]0__2_n_73 ),
        .I1(n_reg[15]),
        .O(\n_reg[2]0_i_18__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_19 
       (.I0(\n_reg[1]0__2_n_88 ),
        .I1(n_reg[0]),
        .O(\n_reg[2]0_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_19__0 
       (.I0(\n_reg[1]0__2_n_74 ),
        .I1(n_reg[14]),
        .O(\n_reg[2]0_i_19__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[2]0_i_1__0 
       (.CI(\n_reg[2]0_i_2__0_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\n_reg[1]0__2_n_61 ,\n_reg[1]0__2_n_62 }),
        .O({\n_reg[2]0_i_1__0_n_4 ,\n_next[1] [31:29]}),
        .S({\<const0>__0__0 ,\n_reg[2]0_i_5__0_n_0 ,\n_reg[2]0_i_6__0_n_0 ,\n_reg[2]0_i_7__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[2]0_i_2 
       (.CI(\n_reg[2]0_i_3_n_0 ),
        .CO({\n_reg[2]0_i_2_n_0 ,\n_reg[2]0_i_2_n_1 ,\n_reg[2]0_i_2_n_2 ,\n_reg[2]0_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[1]0__2_n_79 ,\n_reg[1]0__2_n_80 ,\n_reg[1]0__2_n_81 ,\n_reg[1]0__2_n_82 }),
        .O(\n_next[1] [12:9]),
        .S({\n_reg[2]0_i_10_n_0 ,\n_reg[2]0_i_11_n_0 ,\n_reg[2]0_i_12_n_0 ,\n_reg[2]0_i_13_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_20 
       (.I0(\n_reg[1]0__2_n_89 ),
        .I1(\n_reg[1]0_n_89 ),
        .O(\n_reg[2]0_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_21 
       (.I0(\n_reg[1]0__2_n_90 ),
        .I1(\n_reg[1]0_n_90 ),
        .O(\n_reg[2]0_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[2]0_i_22 
       (.CI(\n_reg[2]0_i_27_n_0 ),
        .CO({\n_reg[2]0_i_22_n_0 ,\n_reg[2]0_i_22_n_1 ,\n_reg[2]0_i_22_n_2 ,\n_reg[2]0_i_22_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[1]0__2_n_95 ,\n_reg[1]0__2_n_96 ,\n_reg[1]0__2_n_97 ,\n_reg[1]0__2_n_98 }),
        .S({\n_reg[2]0_i_28_n_0 ,\n_reg[2]0_i_29_n_0 ,\n_reg[2]0_i_30_n_0 ,\n_reg[2]0_i_31_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_23 
       (.I0(\n_reg[1]0__2_n_91 ),
        .I1(\n_reg[1]0_n_91 ),
        .O(\n_reg[2]0_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_24 
       (.I0(\n_reg[1]0__2_n_92 ),
        .I1(\n_reg[1]0_n_92 ),
        .O(\n_reg[2]0_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_25 
       (.I0(\n_reg[1]0__2_n_93 ),
        .I1(\n_reg[1]0_n_93 ),
        .O(\n_reg[2]0_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_26 
       (.I0(\n_reg[1]0__2_n_94 ),
        .I1(\n_reg[1]0_n_94 ),
        .O(\n_reg[2]0_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[2]0_i_27 
       (.CI(\n_reg[2]0_i_32_n_0 ),
        .CO({\n_reg[2]0_i_27_n_0 ,\n_reg[2]0_i_27_n_1 ,\n_reg[2]0_i_27_n_2 ,\n_reg[2]0_i_27_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[1]0__2_n_99 ,\n_reg[1]0__2_n_100 ,\n_reg[1]0__2_n_101 ,\n_reg[1]0__2_n_102 }),
        .S({\n_reg[2]0_i_33_n_0 ,\n_reg[2]0_i_34_n_0 ,\n_reg[2]0_i_35_n_0 ,\n_reg[2]0_i_36_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_28 
       (.I0(\n_reg[1]0__2_n_95 ),
        .I1(\n_reg[1]0_n_95 ),
        .O(\n_reg[2]0_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_29 
       (.I0(\n_reg[1]0__2_n_96 ),
        .I1(\n_reg[1]0_n_96 ),
        .O(\n_reg[2]0_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[2]0_i_2__0 
       (.CI(\n_reg[2]0_i_3__0_n_0 ),
        .CO({\n_reg[2]0_i_2__0_n_0 ,\n_reg[2]0_i_2__0_n_1 ,\n_reg[2]0_i_2__0_n_2 ,\n_reg[2]0_i_2__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[1]0__2_n_63 ,\n_reg[1]0__2_n_64 ,\n_reg[1]0__2_n_65 ,\n_reg[1]0__2_n_66 }),
        .O(\n_next[1] [28:25]),
        .S({\n_reg[2]0_i_8__0_n_0 ,\n_reg[2]0_i_9__0_n_0 ,\n_reg[2]0_i_10__0_n_0 ,\n_reg[2]0_i_11__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[2]0_i_3 
       (.CI(\n_reg[2]0_i_4_n_0 ),
        .CO({\n_reg[2]0_i_3_n_0 ,\n_reg[2]0_i_3_n_1 ,\n_reg[2]0_i_3_n_2 ,\n_reg[2]0_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[1]0__2_n_83 ,\n_reg[1]0__2_n_84 ,\n_reg[1]0__2_n_85 ,\n_reg[1]0__2_n_86 }),
        .O(\n_next[1] [8:5]),
        .S({\n_reg[2]0_i_14_n_0 ,\n_reg[2]0_i_15_n_0 ,\n_reg[2]0_i_16_n_0 ,\n_reg[2]0_i_17_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_30 
       (.I0(\n_reg[1]0__2_n_97 ),
        .I1(\n_reg[1]0_n_97 ),
        .O(\n_reg[2]0_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_31 
       (.I0(\n_reg[1]0__2_n_98 ),
        .I1(\n_reg[1]0_n_98 ),
        .O(\n_reg[2]0_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[2]0_i_32 
       (.CI(\<const0>__0__0 ),
        .CO({\n_reg[2]0_i_32_n_0 ,\n_reg[2]0_i_32_n_1 ,\n_reg[2]0_i_32_n_2 ,\n_reg[2]0_i_32_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[1]0__2_n_103 ,\n_reg[1]0__2_n_104 ,\n_reg[1]0__2_n_105 ,\<const0>__0__0 }),
        .S({\n_reg[2]0_i_37_n_0 ,\n_reg[2]0_i_38_n_0 ,\n_reg[2]0_i_39_n_0 ,\n_reg[1]0__1_n_89 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_33 
       (.I0(\n_reg[1]0__2_n_99 ),
        .I1(\n_reg[1]0_n_99 ),
        .O(\n_reg[2]0_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_34 
       (.I0(\n_reg[1]0__2_n_100 ),
        .I1(\n_reg[1]0_n_100 ),
        .O(\n_reg[2]0_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_35 
       (.I0(\n_reg[1]0__2_n_101 ),
        .I1(\n_reg[1]0_n_101 ),
        .O(\n_reg[2]0_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_36 
       (.I0(\n_reg[1]0__2_n_102 ),
        .I1(\n_reg[1]0_n_102 ),
        .O(\n_reg[2]0_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_37 
       (.I0(\n_reg[1]0__2_n_103 ),
        .I1(\n_reg[1]0_n_103 ),
        .O(\n_reg[2]0_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_38 
       (.I0(\n_reg[1]0__2_n_104 ),
        .I1(\n_reg[1]0_n_104 ),
        .O(\n_reg[2]0_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_39 
       (.I0(\n_reg[1]0__2_n_105 ),
        .I1(\n_reg[1]0_n_105 ),
        .O(\n_reg[2]0_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[2]0_i_3__0 
       (.CI(\n_reg[2]0_i_4__0_n_0 ),
        .CO({\n_reg[2]0_i_3__0_n_0 ,\n_reg[2]0_i_3__0_n_1 ,\n_reg[2]0_i_3__0_n_2 ,\n_reg[2]0_i_3__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[1]0__2_n_67 ,\n_reg[1]0__2_n_68 ,\n_reg[1]0__2_n_69 ,\n_reg[1]0__2_n_70 }),
        .O(\n_next[1] [24:21]),
        .S({\n_reg[2]0_i_12__0_n_0 ,\n_reg[2]0_i_13__0_n_0 ,\n_reg[2]0_i_14__0_n_0 ,\n_reg[2]0_i_15__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[2]0_i_4 
       (.CI(\n_reg[2]0_i_5_n_0 ),
        .CO({\n_reg[2]0_i_4_n_0 ,\n_reg[2]0_i_4_n_1 ,\n_reg[2]0_i_4_n_2 ,\n_reg[2]0_i_4_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[1]0__2_n_87 ,\n_reg[1]0__2_n_88 ,\n_reg[1]0__2_n_89 ,\n_reg[1]0__2_n_90 }),
        .O(\n_next[1] [4:1]),
        .S({\n_reg[2]0_i_18_n_0 ,\n_reg[2]0_i_19_n_0 ,\n_reg[2]0_i_20_n_0 ,\n_reg[2]0_i_21_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[2]0_i_4__0 
       (.CI(\n_reg[2]0_i_1_n_0 ),
        .CO({\n_reg[2]0_i_4__0_n_0 ,\n_reg[2]0_i_4__0_n_1 ,\n_reg[2]0_i_4__0_n_2 ,\n_reg[2]0_i_4__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[1]0__2_n_71 ,\n_reg[1]0__2_n_72 ,\n_reg[1]0__2_n_73 ,\n_reg[1]0__2_n_74 }),
        .O(\n_next[1] [20:17]),
        .S({\n_reg[2]0_i_16__0_n_0 ,\n_reg[2]0_i_17__0_n_0 ,\n_reg[2]0_i_18__0_n_0 ,\n_reg[2]0_i_19__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[2]0_i_5 
       (.CI(\n_reg[2]0_i_22_n_0 ),
        .CO({\n_reg[2]0_i_5_n_0 ,\n_reg[2]0_i_5_n_1 ,\n_reg[2]0_i_5_n_2 ,\n_reg[2]0_i_5_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[1]0__2_n_91 ,\n_reg[1]0__2_n_92 ,\n_reg[1]0__2_n_93 ,\n_reg[1]0__2_n_94 }),
        .O({\n_next[1] [0],\n_reg[2]0_i_5_n_5 ,\n_reg[2]0_i_5_n_6 ,\n_reg[2]0_i_5_n_7 }),
        .S({\n_reg[2]0_i_23_n_0 ,\n_reg[2]0_i_24_n_0 ,\n_reg[2]0_i_25_n_0 ,\n_reg[2]0_i_26_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_5__0 
       (.I0(\n_reg[1]0__2_n_60 ),
        .I1(n_reg[28]),
        .O(\n_reg[2]0_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_6 
       (.I0(\n_reg[1]0__2_n_75 ),
        .I1(n_reg[13]),
        .O(\n_reg[2]0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_6__0 
       (.I0(\n_reg[1]0__2_n_61 ),
        .I1(n_reg[27]),
        .O(\n_reg[2]0_i_6__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_7 
       (.I0(\n_reg[1]0__2_n_76 ),
        .I1(n_reg[12]),
        .O(\n_reg[2]0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_7__0 
       (.I0(\n_reg[1]0__2_n_62 ),
        .I1(n_reg[26]),
        .O(\n_reg[2]0_i_7__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_8 
       (.I0(\n_reg[1]0__2_n_77 ),
        .I1(n_reg[11]),
        .O(\n_reg[2]0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_8__0 
       (.I0(\n_reg[1]0__2_n_63 ),
        .I1(n_reg[25]),
        .O(\n_reg[2]0_i_8__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_9 
       (.I0(\n_reg[1]0__2_n_78 ),
        .I1(n_reg[10]),
        .O(\n_reg[2]0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[2]0_i_9__0 
       (.I0(\n_reg[1]0__2_n_64 ),
        .I1(n_reg[24]),
        .O(\n_reg[2]0_i_9__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-10 {cell *THIS*} {string 16x18 4}}" *) 
  DSP48E1 #(
    .ACASCREG(1),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(1),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(1),
    .BREG(1),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \n_reg[3]0 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\r_reg[2]0 [16:1],\n_reg[3]0_i_9__1_n_7 }),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\n_next[2] [31:17]}),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const1>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const1>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\n_reg[3]0_n_58 ,\n_reg[3]0_n_59 ,\n_reg[3]0_n_60 ,\n_reg[3]0_n_61 ,\n_reg[3]0_n_62 ,\n_reg[3]0_n_63 ,\n_reg[3]0_n_64 ,\n_reg[3]0_n_65 ,\n_reg[3]0_n_66 ,\n_reg[3]0_n_67 ,\n_reg[3]0_n_68 ,\n_reg[3]0_n_69 ,\n_reg[3]0_n_70 ,\n_reg[3]0_n_71 ,\n_reg[3]0_n_72 ,\n_reg[3]0_n_73 ,\n_reg[3]0_n_74 ,\n_reg[3]0_n_75 ,\n_reg[3]0_n_76 ,\n_reg[3]0_n_77 ,\n_reg[3]0_n_78 ,\n_reg[3]0_n_79 ,\n_reg[3]0_n_80 ,\n_reg[3]0_n_81 ,\n_reg[3]0_n_82 ,\n_reg[3]0_n_83 ,\n_reg[3]0_n_84 ,\n_reg[3]0_n_85 ,\n_reg[3]0_n_86 ,\n_reg[3]0_n_87 ,\n_reg[3]0_n_88 ,\n_reg[3]0_n_89 ,\n_reg[3]0_n_90 ,\n_reg[3]0_n_91 ,\n_reg[3]0_n_92 ,\n_reg[3]0_n_93 ,\n_reg[3]0_n_94 ,\n_reg[3]0_n_95 ,\n_reg[3]0_n_96 ,\n_reg[3]0_n_97 ,\n_reg[3]0_n_98 ,\n_reg[3]0_n_99 ,\n_reg[3]0_n_100 ,\n_reg[3]0_n_101 ,\n_reg[3]0_n_102 ,\n_reg[3]0_n_103 ,\n_reg[3]0_n_104 ,\n_reg[3]0_n_105 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .PCOUT({\n_reg[3]0_n_106 ,\n_reg[3]0_n_107 ,\n_reg[3]0_n_108 ,\n_reg[3]0_n_109 ,\n_reg[3]0_n_110 ,\n_reg[3]0_n_111 ,\n_reg[3]0_n_112 ,\n_reg[3]0_n_113 ,\n_reg[3]0_n_114 ,\n_reg[3]0_n_115 ,\n_reg[3]0_n_116 ,\n_reg[3]0_n_117 ,\n_reg[3]0_n_118 ,\n_reg[3]0_n_119 ,\n_reg[3]0_n_120 ,\n_reg[3]0_n_121 ,\n_reg[3]0_n_122 ,\n_reg[3]0_n_123 ,\n_reg[3]0_n_124 ,\n_reg[3]0_n_125 ,\n_reg[3]0_n_126 ,\n_reg[3]0_n_127 ,\n_reg[3]0_n_128 ,\n_reg[3]0_n_129 ,\n_reg[3]0_n_130 ,\n_reg[3]0_n_131 ,\n_reg[3]0_n_132 ,\n_reg[3]0_n_133 ,\n_reg[3]0_n_134 ,\n_reg[3]0_n_135 ,\n_reg[3]0_n_136 ,\n_reg[3]0_n_137 ,\n_reg[3]0_n_138 ,\n_reg[3]0_n_139 ,\n_reg[3]0_n_140 ,\n_reg[3]0_n_141 ,\n_reg[3]0_n_142 ,\n_reg[3]0_n_143 ,\n_reg[3]0_n_144 ,\n_reg[3]0_n_145 ,\n_reg[3]0_n_146 ,\n_reg[3]0_n_147 ,\n_reg[3]0_n_148 ,\n_reg[3]0_n_149 ,\n_reg[3]0_n_150 ,\n_reg[3]0_n_151 ,\n_reg[3]0_n_152 ,\n_reg[3]0_n_153 }),
        .RSTA(RSTA),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(RSTA),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-10 {cell *THIS*} {string 16x16 4}}" *) 
  DSP48E1 #(
    .ACASCREG(1),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(1),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(1),
    .BREG(1),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \n_reg[3]0__0 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\n_next[2] [31:17]}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\r_reg[2]0 [31:17]}),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const1>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const1>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\n_reg[3]0__0_n_58 ,\n_reg[3]0__0_n_59 ,\n_reg[3]0__0_n_60 ,\n_reg[3]0__0_n_61 ,\n_reg[3]0__0_n_62 ,\n_reg[3]0__0_n_63 ,\n_reg[3]0__0_n_64 ,\n_reg[3]0__0_n_65 ,\n_reg[3]0__0_n_66 ,\n_reg[3]0__0_n_67 ,\n_reg[3]0__0_n_68 ,\n_reg[3]0__0_n_69 ,\n_reg[3]0__0_n_70 ,\n_reg[3]0__0_n_71 ,\n_reg[3]0__0_n_72 ,\n_reg[3]0__0_n_73 ,\n_reg[3]0__0_n_74 ,\n_reg[3]0__0_n_75 ,\n_reg[3]0__0_n_76 ,\n_reg[3]0__0_n_77 ,\n_reg[3]0__0_n_78 ,\n_reg[3]0__0_n_79 ,\n_reg[3]0__0_n_80 ,\n_reg[3]0__0_n_81 ,\n_reg[3]0__0_n_82 ,\n_reg[3]0__0_n_83 ,\n_reg[3]0__0_n_84 ,\n_reg[3]0__0_n_85 ,\n_reg[3]0__0_n_86 ,\n_reg[3]0__0_n_87 ,\n_reg[3]0__0_n_88 ,\n_reg[3]0__0_n_89 ,\n_reg[3]0__0_n_90 ,\n_reg[3]0__0_n_91 ,\n_reg[3]0__0_n_92 ,\n_reg[3]0__0_n_93 ,\n_reg[3]0__0_n_94 ,\n_reg[3]0__0_n_95 ,\n_reg[3]0__0_n_96 ,\n_reg[3]0__0_n_97 ,\n_reg[3]0__0_n_98 ,\n_reg[3]0__0_n_99 ,\n_reg[3]0__0_n_100 ,\n_reg[3]0__0_n_101 ,\n_reg[3]0__0_n_102 ,\n_reg[3]0__0_n_103 ,\n_reg[3]0__0_n_104 ,\n_reg[3]0__0_n_105 }),
        .PCIN({\n_reg[3]0_n_106 ,\n_reg[3]0_n_107 ,\n_reg[3]0_n_108 ,\n_reg[3]0_n_109 ,\n_reg[3]0_n_110 ,\n_reg[3]0_n_111 ,\n_reg[3]0_n_112 ,\n_reg[3]0_n_113 ,\n_reg[3]0_n_114 ,\n_reg[3]0_n_115 ,\n_reg[3]0_n_116 ,\n_reg[3]0_n_117 ,\n_reg[3]0_n_118 ,\n_reg[3]0_n_119 ,\n_reg[3]0_n_120 ,\n_reg[3]0_n_121 ,\n_reg[3]0_n_122 ,\n_reg[3]0_n_123 ,\n_reg[3]0_n_124 ,\n_reg[3]0_n_125 ,\n_reg[3]0_n_126 ,\n_reg[3]0_n_127 ,\n_reg[3]0_n_128 ,\n_reg[3]0_n_129 ,\n_reg[3]0_n_130 ,\n_reg[3]0_n_131 ,\n_reg[3]0_n_132 ,\n_reg[3]0_n_133 ,\n_reg[3]0_n_134 ,\n_reg[3]0_n_135 ,\n_reg[3]0_n_136 ,\n_reg[3]0_n_137 ,\n_reg[3]0_n_138 ,\n_reg[3]0_n_139 ,\n_reg[3]0_n_140 ,\n_reg[3]0_n_141 ,\n_reg[3]0_n_142 ,\n_reg[3]0_n_143 ,\n_reg[3]0_n_144 ,\n_reg[3]0_n_145 ,\n_reg[3]0_n_146 ,\n_reg[3]0_n_147 ,\n_reg[3]0_n_148 ,\n_reg[3]0_n_149 ,\n_reg[3]0_n_150 ,\n_reg[3]0_n_151 ,\n_reg[3]0_n_152 ,\n_reg[3]0_n_153 }),
        .RSTA(RSTA),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(RSTA),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-10 {cell *THIS*} {string 18x18 4}}" *) 
  DSP48E1 #(
    .ACASCREG(1),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(1),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(1),
    .BREG(1),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \n_reg[3]0__1 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\n_next[2] [16:0]}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ACOUT({\n_reg[3]0__1_n_24 ,\n_reg[3]0__1_n_25 ,\n_reg[3]0__1_n_26 ,\n_reg[3]0__1_n_27 ,\n_reg[3]0__1_n_28 ,\n_reg[3]0__1_n_29 ,\n_reg[3]0__1_n_30 ,\n_reg[3]0__1_n_31 ,\n_reg[3]0__1_n_32 ,\n_reg[3]0__1_n_33 ,\n_reg[3]0__1_n_34 ,\n_reg[3]0__1_n_35 ,\n_reg[3]0__1_n_36 ,\n_reg[3]0__1_n_37 ,\n_reg[3]0__1_n_38 ,\n_reg[3]0__1_n_39 ,\n_reg[3]0__1_n_40 ,\n_reg[3]0__1_n_41 ,\n_reg[3]0__1_n_42 ,\n_reg[3]0__1_n_43 ,\n_reg[3]0__1_n_44 ,\n_reg[3]0__1_n_45 ,\n_reg[3]0__1_n_46 ,\n_reg[3]0__1_n_47 ,\n_reg[3]0__1_n_48 ,\n_reg[3]0__1_n_49 ,\n_reg[3]0__1_n_50 ,\n_reg[3]0__1_n_51 ,\n_reg[3]0__1_n_52 ,\n_reg[3]0__1_n_53 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\r_reg[2]0 [16:1],\n_reg[3]0_i_9__1_n_7 }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const1>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const1>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\n_reg[3]0__1_n_58 ,\n_reg[3]0__1_n_59 ,\n_reg[3]0__1_n_60 ,\n_reg[3]0__1_n_61 ,\n_reg[3]0__1_n_62 ,\n_reg[3]0__1_n_63 ,\n_reg[3]0__1_n_64 ,\n_reg[3]0__1_n_65 ,\n_reg[3]0__1_n_66 ,\n_reg[3]0__1_n_67 ,\n_reg[3]0__1_n_68 ,\n_reg[3]0__1_n_69 ,\n_reg[3]0__1_n_70 ,\n_reg[3]0__1_n_71 ,\n_reg[3]0__1_n_72 ,\n_reg[3]0__1_n_73 ,\n_reg[3]0__1_n_74 ,\n_reg[3]0__1_n_75 ,\n_reg[3]0__1_n_76 ,\n_reg[3]0__1_n_77 ,\n_reg[3]0__1_n_78 ,\n_reg[3]0__1_n_79 ,\n_reg[3]0__1_n_80 ,\n_reg[3]0__1_n_81 ,\n_reg[3]0__1_n_82 ,\n_reg[3]0__1_n_83 ,\n_reg[3]0__1_n_84 ,\n_reg[3]0__1_n_85 ,\n_reg[3]0__1_n_86 ,\n_reg[3]0__1_n_87 ,\n_reg[3]0__1_n_88 ,\n_reg[3]0__1_n_89 ,\n_reg[3]0__1_n_90 ,\n_reg[3]0__1_n_91 ,\n_reg[3]0__1_n_92 ,\n_reg[3]0__1_n_93 ,\n_reg[3]0__1_n_94 ,\n_reg[3]0__1_n_95 ,\n_reg[3]0__1_n_96 ,\n_reg[3]0__1_n_97 ,\n_reg[3]0__1_n_98 ,\n_reg[3]0__1_n_99 ,\n_reg[3]0__1_n_100 ,\n_reg[3]0__1_n_101 ,\n_reg[3]0__1_n_102 ,\n_reg[3]0__1_n_103 ,\n_reg[3]0__1_n_104 ,\n_reg[3]0__1_n_105 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .PCOUT({\n_reg[3]0__1_n_106 ,\n_reg[3]0__1_n_107 ,\n_reg[3]0__1_n_108 ,\n_reg[3]0__1_n_109 ,\n_reg[3]0__1_n_110 ,\n_reg[3]0__1_n_111 ,\n_reg[3]0__1_n_112 ,\n_reg[3]0__1_n_113 ,\n_reg[3]0__1_n_114 ,\n_reg[3]0__1_n_115 ,\n_reg[3]0__1_n_116 ,\n_reg[3]0__1_n_117 ,\n_reg[3]0__1_n_118 ,\n_reg[3]0__1_n_119 ,\n_reg[3]0__1_n_120 ,\n_reg[3]0__1_n_121 ,\n_reg[3]0__1_n_122 ,\n_reg[3]0__1_n_123 ,\n_reg[3]0__1_n_124 ,\n_reg[3]0__1_n_125 ,\n_reg[3]0__1_n_126 ,\n_reg[3]0__1_n_127 ,\n_reg[3]0__1_n_128 ,\n_reg[3]0__1_n_129 ,\n_reg[3]0__1_n_130 ,\n_reg[3]0__1_n_131 ,\n_reg[3]0__1_n_132 ,\n_reg[3]0__1_n_133 ,\n_reg[3]0__1_n_134 ,\n_reg[3]0__1_n_135 ,\n_reg[3]0__1_n_136 ,\n_reg[3]0__1_n_137 ,\n_reg[3]0__1_n_138 ,\n_reg[3]0__1_n_139 ,\n_reg[3]0__1_n_140 ,\n_reg[3]0__1_n_141 ,\n_reg[3]0__1_n_142 ,\n_reg[3]0__1_n_143 ,\n_reg[3]0__1_n_144 ,\n_reg[3]0__1_n_145 ,\n_reg[3]0__1_n_146 ,\n_reg[3]0__1_n_147 ,\n_reg[3]0__1_n_148 ,\n_reg[3]0__1_n_149 ,\n_reg[3]0__1_n_150 ,\n_reg[3]0__1_n_151 ,\n_reg[3]0__1_n_152 ,\n_reg[3]0__1_n_153 }),
        .RSTA(RSTA),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(RSTA),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-10 {cell *THIS*} {string 18x16 4}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("CASCADE"),
    .BCASCREG(1),
    .BREG(1),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \n_reg[3]0__2 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ACIN({\n_reg[3]0__1_n_24 ,\n_reg[3]0__1_n_25 ,\n_reg[3]0__1_n_26 ,\n_reg[3]0__1_n_27 ,\n_reg[3]0__1_n_28 ,\n_reg[3]0__1_n_29 ,\n_reg[3]0__1_n_30 ,\n_reg[3]0__1_n_31 ,\n_reg[3]0__1_n_32 ,\n_reg[3]0__1_n_33 ,\n_reg[3]0__1_n_34 ,\n_reg[3]0__1_n_35 ,\n_reg[3]0__1_n_36 ,\n_reg[3]0__1_n_37 ,\n_reg[3]0__1_n_38 ,\n_reg[3]0__1_n_39 ,\n_reg[3]0__1_n_40 ,\n_reg[3]0__1_n_41 ,\n_reg[3]0__1_n_42 ,\n_reg[3]0__1_n_43 ,\n_reg[3]0__1_n_44 ,\n_reg[3]0__1_n_45 ,\n_reg[3]0__1_n_46 ,\n_reg[3]0__1_n_47 ,\n_reg[3]0__1_n_48 ,\n_reg[3]0__1_n_49 ,\n_reg[3]0__1_n_50 ,\n_reg[3]0__1_n_51 ,\n_reg[3]0__1_n_52 ,\n_reg[3]0__1_n_53 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\r_reg[2]0 [31:17]}),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const1>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\n_reg[3]0__2_n_58 ,\n_reg[3]0__2_n_59 ,\n_reg[3]0__2_n_60 ,\n_reg[3]0__2_n_61 ,\n_reg[3]0__2_n_62 ,\n_reg[3]0__2_n_63 ,\n_reg[3]0__2_n_64 ,\n_reg[3]0__2_n_65 ,\n_reg[3]0__2_n_66 ,\n_reg[3]0__2_n_67 ,\n_reg[3]0__2_n_68 ,\n_reg[3]0__2_n_69 ,\n_reg[3]0__2_n_70 ,\n_reg[3]0__2_n_71 ,\n_reg[3]0__2_n_72 ,\n_reg[3]0__2_n_73 ,\n_reg[3]0__2_n_74 ,\n_reg[3]0__2_n_75 ,\n_reg[3]0__2_n_76 ,\n_reg[3]0__2_n_77 ,\n_reg[3]0__2_n_78 ,\n_reg[3]0__2_n_79 ,\n_reg[3]0__2_n_80 ,\n_reg[3]0__2_n_81 ,\n_reg[3]0__2_n_82 ,\n_reg[3]0__2_n_83 ,\n_reg[3]0__2_n_84 ,\n_reg[3]0__2_n_85 ,\n_reg[3]0__2_n_86 ,\n_reg[3]0__2_n_87 ,\n_reg[3]0__2_n_88 ,\n_reg[3]0__2_n_89 ,\n_reg[3]0__2_n_90 ,\n_reg[3]0__2_n_91 ,\n_reg[3]0__2_n_92 ,\n_reg[3]0__2_n_93 ,\n_reg[3]0__2_n_94 ,\n_reg[3]0__2_n_95 ,\n_reg[3]0__2_n_96 ,\n_reg[3]0__2_n_97 ,\n_reg[3]0__2_n_98 ,\n_reg[3]0__2_n_99 ,\n_reg[3]0__2_n_100 ,\n_reg[3]0__2_n_101 ,\n_reg[3]0__2_n_102 ,\n_reg[3]0__2_n_103 ,\n_reg[3]0__2_n_104 ,\n_reg[3]0__2_n_105 }),
        .PCIN({\n_reg[3]0__1_n_106 ,\n_reg[3]0__1_n_107 ,\n_reg[3]0__1_n_108 ,\n_reg[3]0__1_n_109 ,\n_reg[3]0__1_n_110 ,\n_reg[3]0__1_n_111 ,\n_reg[3]0__1_n_112 ,\n_reg[3]0__1_n_113 ,\n_reg[3]0__1_n_114 ,\n_reg[3]0__1_n_115 ,\n_reg[3]0__1_n_116 ,\n_reg[3]0__1_n_117 ,\n_reg[3]0__1_n_118 ,\n_reg[3]0__1_n_119 ,\n_reg[3]0__1_n_120 ,\n_reg[3]0__1_n_121 ,\n_reg[3]0__1_n_122 ,\n_reg[3]0__1_n_123 ,\n_reg[3]0__1_n_124 ,\n_reg[3]0__1_n_125 ,\n_reg[3]0__1_n_126 ,\n_reg[3]0__1_n_127 ,\n_reg[3]0__1_n_128 ,\n_reg[3]0__1_n_129 ,\n_reg[3]0__1_n_130 ,\n_reg[3]0__1_n_131 ,\n_reg[3]0__1_n_132 ,\n_reg[3]0__1_n_133 ,\n_reg[3]0__1_n_134 ,\n_reg[3]0__1_n_135 ,\n_reg[3]0__1_n_136 ,\n_reg[3]0__1_n_137 ,\n_reg[3]0__1_n_138 ,\n_reg[3]0__1_n_139 ,\n_reg[3]0__1_n_140 ,\n_reg[3]0__1_n_141 ,\n_reg[3]0__1_n_142 ,\n_reg[3]0__1_n_143 ,\n_reg[3]0__1_n_144 ,\n_reg[3]0__1_n_145 ,\n_reg[3]0__1_n_146 ,\n_reg[3]0__1_n_147 ,\n_reg[3]0__1_n_148 ,\n_reg[3]0__1_n_149 ,\n_reg[3]0__1_n_150 ,\n_reg[3]0__1_n_151 ,\n_reg[3]0__1_n_152 ,\n_reg[3]0__1_n_153 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(RSTA),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_1 
       (.CI(\n_reg[3]0_i_2_n_0 ),
        .CO({\n_reg[3]0_i_1_n_0 ,\n_reg[3]0_i_1_n_1 ,\n_reg[3]0_i_1_n_2 ,\n_reg[3]0_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[2]0__2_n_75 ,\n_reg[2]0__2_n_76 ,\n_reg[2]0__2_n_77 ,\n_reg[2]0__2_n_78 }),
        .O(\n_next[2] [16:13]),
        .S({\n_reg[3]0_i_6_n_0 ,\n_reg[3]0_i_7_n_0 ,\n_reg[3]0_i_8_n_0 ,\n_reg[3]0_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_10 
       (.I0(\n_reg[2]0__2_n_79 ),
        .I1(\n_reg[2]0__0_n_96 ),
        .O(\n_reg[3]0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_10__0 
       (.I0(\n_reg[2]0__2_n_60 ),
        .I1(\n_reg[2]0__0_n_77 ),
        .O(\n_reg[3]0_i_10__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_10__1 
       (.I0(\n_reg[3]0_i_21__1_n_5 ),
        .O(\n_reg[3]0_i_10__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_11 
       (.I0(\n_reg[2]0__2_n_80 ),
        .I1(\n_reg[2]0__0_n_97 ),
        .O(\n_reg[3]0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_11__0 
       (.I0(\n_reg[2]0__2_n_61 ),
        .I1(\n_reg[2]0__0_n_78 ),
        .O(\n_reg[3]0_i_11__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_11__1 
       (.I0(\n_reg[3]0_i_21__1_n_6 ),
        .O(\n_reg[3]0_i_11__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_12 
       (.I0(\n_reg[2]0__2_n_81 ),
        .I1(\n_reg[2]0__0_n_98 ),
        .O(\n_reg[3]0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_12__0 
       (.I0(\n_reg[2]0__2_n_62 ),
        .I1(\n_reg[2]0__0_n_79 ),
        .O(\n_reg[3]0_i_12__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_12__1 
       (.I0(\n_reg[3]0_i_21__1_n_7 ),
        .O(\n_reg[3]0_i_12__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_13 
       (.I0(\n_reg[2]0__2_n_82 ),
        .I1(\n_reg[2]0__0_n_99 ),
        .O(\n_reg[3]0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_13__0 
       (.I0(\n_reg[2]0__2_n_63 ),
        .I1(\n_reg[2]0__0_n_80 ),
        .O(\n_reg[3]0_i_13__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_13__1 
       (.I0(\n_reg[3]0_i_22__1_n_4 ),
        .O(\n_reg[3]0_i_13__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_14 
       (.I0(\n_reg[2]0__2_n_83 ),
        .I1(\n_reg[2]0__0_n_100 ),
        .O(\n_reg[3]0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_14__0 
       (.I0(\n_reg[2]0__2_n_64 ),
        .I1(\n_reg[2]0__0_n_81 ),
        .O(\n_reg[3]0_i_14__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_14__1 
       (.I0(\n_reg[3]0_i_22__1_n_5 ),
        .O(\n_reg[3]0_i_14__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_15 
       (.I0(\n_reg[2]0__2_n_84 ),
        .I1(\n_reg[2]0__0_n_101 ),
        .O(\n_reg[3]0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_15__0 
       (.I0(\n_reg[2]0__2_n_65 ),
        .I1(\n_reg[2]0__0_n_82 ),
        .O(\n_reg[3]0_i_15__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_15__1 
       (.I0(\n_reg[3]0_i_22__1_n_6 ),
        .O(\n_reg[3]0_i_15__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_16 
       (.I0(\n_reg[2]0__2_n_85 ),
        .I1(\n_reg[2]0__0_n_102 ),
        .O(\n_reg[3]0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_16__0 
       (.I0(\n_reg[2]0__2_n_66 ),
        .I1(\n_reg[2]0__0_n_83 ),
        .O(\n_reg[3]0_i_16__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_16__1 
       (.I0(\n_reg[3]0_i_22__1_n_7 ),
        .O(\n_reg[3]0_i_16__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_17 
       (.I0(\n_reg[2]0__2_n_86 ),
        .I1(\n_reg[2]0__0_n_103 ),
        .O(\n_reg[3]0_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_17__0 
       (.I0(\n_reg[2]0__2_n_67 ),
        .I1(\n_reg[2]0__0_n_84 ),
        .O(\n_reg[3]0_i_17__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_17__1 
       (.I0(\n_reg[3]0_i_47_n_4 ),
        .O(\n_reg[3]0_i_17__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_18 
       (.I0(\n_reg[2]0__2_n_87 ),
        .I1(\n_reg[2]0__0_n_104 ),
        .O(\n_reg[3]0_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_18__0 
       (.I0(\n_reg[2]0__2_n_68 ),
        .I1(\n_reg[2]0__0_n_85 ),
        .O(\n_reg[3]0_i_18__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_18__1 
       (.I0(\n_reg[3]0_i_47_n_5 ),
        .O(\n_reg[3]0_i_18__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_19 
       (.I0(\n_reg[2]0__2_n_88 ),
        .I1(\n_reg[2]0__0_n_105 ),
        .O(\n_reg[3]0_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_19__0 
       (.I0(\n_reg[2]0__2_n_69 ),
        .I1(\n_reg[2]0__0_n_86 ),
        .O(\n_reg[3]0_i_19__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_19__1 
       (.I0(\n_reg[3]0_i_47_n_6 ),
        .O(\n_reg[3]0_i_19__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_1__0 
       (.CI(\n_reg[3]0_i_2__0_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\n_reg[2]0__2_n_61 ,\n_reg[2]0__2_n_62 }),
        .O({\n_reg[3]0_i_1__0_n_4 ,\n_next[2] [31:29]}),
        .S({\<const0>__0__0 ,\n_reg[3]0_i_10__0_n_0 ,\n_reg[3]0_i_11__0_n_0 ,\n_reg[3]0_i_12__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_1__1 
       (.CI(\n_reg[3]0_i_2__1_n_0 ),
        .CO({\n_reg[3]0_i_1__1_n_0 ,\r_reg[2]0 [31],\n_reg[3]0_i_1__1_n_2 ,\n_reg[3]0_i_1__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\n_reg[3]0_i_5__0_n_0 ,\<const0>__0__0 }),
        .O({\n_reg[3]0_i_1__1_n_4 ,\n_reg[3]0_i_1__1_n_5 ,\r_reg[2]0 [30:29]}),
        .S({\<const0>__0__0 ,\<const1>__0__0 ,\n_reg[3]0_i_20__1_n_5 ,\n_reg[3]0_i_7__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_2 
       (.CI(\n_reg[3]0_i_3_n_0 ),
        .CO({\n_reg[3]0_i_2_n_0 ,\n_reg[3]0_i_2_n_1 ,\n_reg[3]0_i_2_n_2 ,\n_reg[3]0_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[2]0__2_n_79 ,\n_reg[2]0__2_n_80 ,\n_reg[2]0__2_n_81 ,\n_reg[2]0__2_n_82 }),
        .O(\n_next[2] [12:9]),
        .S({\n_reg[3]0_i_10_n_0 ,\n_reg[3]0_i_11_n_0 ,\n_reg[3]0_i_12_n_0 ,\n_reg[3]0_i_13_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_20 
       (.I0(\n_reg[2]0__2_n_89 ),
        .I1(\n_reg[2]0_n_89 ),
        .O(\n_reg[3]0_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_20__0 
       (.I0(\n_reg[2]0__2_n_70 ),
        .I1(\n_reg[2]0__0_n_87 ),
        .O(\n_reg[3]0_i_20__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_20__1 
       (.CI(\n_reg[3]0_i_21__1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\r_reg[2]1__2_n_61 ,\r_reg[2]1__2_n_62 }),
        .O({\n_reg[3]0_i_20__1_n_4 ,\n_reg[3]0_i_20__1_n_5 ,\n_reg[3]0_i_20__1_n_6 ,\n_reg[3]0_i_20__1_n_7 }),
        .S({\<const0>__0__0 ,\n_reg[3]0_i_23__1_n_0 ,\n_reg[3]0_i_24__1_n_0 ,\n_reg[3]0_i_25__1_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_21 
       (.I0(\n_reg[2]0__2_n_90 ),
        .I1(\n_reg[2]0_n_90 ),
        .O(\n_reg[3]0_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_21__0 
       (.I0(\n_reg[2]0__2_n_71 ),
        .I1(\n_reg[2]0__0_n_88 ),
        .O(\n_reg[3]0_i_21__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_21__1 
       (.CI(\n_reg[3]0_i_22__1_n_0 ),
        .CO({\n_reg[3]0_i_21__1_n_0 ,\n_reg[3]0_i_21__1_n_1 ,\n_reg[3]0_i_21__1_n_2 ,\n_reg[3]0_i_21__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\r_reg[2]1__2_n_63 ,\r_reg[2]1__2_n_64 ,\r_reg[2]1__2_n_65 ,\r_reg[2]1__2_n_66 }),
        .O({\n_reg[3]0_i_21__1_n_4 ,\n_reg[3]0_i_21__1_n_5 ,\n_reg[3]0_i_21__1_n_6 ,\n_reg[3]0_i_21__1_n_7 }),
        .S({\n_reg[3]0_i_26__1_n_0 ,\n_reg[3]0_i_27__1_n_0 ,\n_reg[3]0_i_28__1_n_0 ,\n_reg[3]0_i_29__1_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_22 
       (.CI(\n_reg[3]0_i_27_n_0 ),
        .CO({\n_reg[3]0_i_22_n_0 ,\n_reg[3]0_i_22_n_1 ,\n_reg[3]0_i_22_n_2 ,\n_reg[3]0_i_22_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[2]0__2_n_95 ,\n_reg[2]0__2_n_96 ,\n_reg[2]0__2_n_97 ,\n_reg[2]0__2_n_98 }),
        .S({\n_reg[3]0_i_28_n_0 ,\n_reg[3]0_i_29_n_0 ,\n_reg[3]0_i_30_n_0 ,\n_reg[3]0_i_31_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_22__0 
       (.I0(\n_reg[2]0__2_n_72 ),
        .I1(\n_reg[2]0__0_n_89 ),
        .O(\n_reg[3]0_i_22__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_22__1 
       (.CI(\n_reg[3]0_i_47_n_0 ),
        .CO({\n_reg[3]0_i_22__1_n_0 ,\n_reg[3]0_i_22__1_n_1 ,\n_reg[3]0_i_22__1_n_2 ,\n_reg[3]0_i_22__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\r_reg[2]1__2_n_67 ,\r_reg[2]1__2_n_68 ,\r_reg[2]1__2_n_69 ,\r_reg[2]1__2_n_70 }),
        .O({\n_reg[3]0_i_22__1_n_4 ,\n_reg[3]0_i_22__1_n_5 ,\n_reg[3]0_i_22__1_n_6 ,\n_reg[3]0_i_22__1_n_7 }),
        .S({\n_reg[3]0_i_30__1_n_0 ,\n_reg[3]0_i_31__1_n_0 ,\n_reg[3]0_i_32__1_n_0 ,\n_reg[3]0_i_33__1_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_23 
       (.I0(\n_reg[2]0__2_n_91 ),
        .I1(\n_reg[2]0_n_91 ),
        .O(\n_reg[3]0_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_23__0 
       (.I0(\n_reg[2]0__2_n_73 ),
        .I1(\n_reg[2]0__0_n_90 ),
        .O(\n_reg[3]0_i_23__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_23__1 
       (.I0(\r_reg[2]1__2_n_60 ),
        .I1(r_reg[28]),
        .O(\n_reg[3]0_i_23__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_24 
       (.I0(\n_reg[2]0__2_n_92 ),
        .I1(\n_reg[2]0_n_92 ),
        .O(\n_reg[3]0_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_24__0 
       (.I0(\n_reg[2]0__2_n_74 ),
        .I1(\n_reg[2]0__0_n_91 ),
        .O(\n_reg[3]0_i_24__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_24__1 
       (.I0(\r_reg[2]1__2_n_61 ),
        .I1(r_reg[27]),
        .O(\n_reg[3]0_i_24__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_25 
       (.I0(\n_reg[2]0__2_n_93 ),
        .I1(\n_reg[2]0_n_93 ),
        .O(\n_reg[3]0_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_25__0 
       (.I0(\n_reg[3]0_i_47_n_7 ),
        .O(\n_reg[3]0_i_25__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_25__1 
       (.I0(\r_reg[2]1__2_n_62 ),
        .I1(r_reg[26]),
        .O(\n_reg[3]0_i_25__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_26 
       (.I0(\n_reg[2]0__2_n_94 ),
        .I1(\n_reg[2]0_n_94 ),
        .O(\n_reg[3]0_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_26__0 
       (.I0(\n_reg[3]0_i_48_n_4 ),
        .O(\n_reg[3]0_i_26__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_26__1 
       (.I0(\r_reg[2]1__2_n_63 ),
        .I1(r_reg[25]),
        .O(\n_reg[3]0_i_26__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_27 
       (.CI(\n_reg[3]0_i_32_n_0 ),
        .CO({\n_reg[3]0_i_27_n_0 ,\n_reg[3]0_i_27_n_1 ,\n_reg[3]0_i_27_n_2 ,\n_reg[3]0_i_27_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[2]0__2_n_99 ,\n_reg[2]0__2_n_100 ,\n_reg[2]0__2_n_101 ,\n_reg[2]0__2_n_102 }),
        .S({\n_reg[3]0_i_33_n_0 ,\n_reg[3]0_i_34_n_0 ,\n_reg[3]0_i_35_n_0 ,\n_reg[3]0_i_36_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_27__0 
       (.I0(\n_reg[3]0_i_48_n_5 ),
        .O(\n_reg[3]0_i_27__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_27__1 
       (.I0(\r_reg[2]1__2_n_64 ),
        .I1(r_reg[24]),
        .O(\n_reg[3]0_i_27__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_28 
       (.I0(\n_reg[2]0__2_n_95 ),
        .I1(\n_reg[2]0_n_95 ),
        .O(\n_reg[3]0_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_28__0 
       (.I0(\n_reg[3]0_i_48_n_6 ),
        .O(\n_reg[3]0_i_28__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_28__1 
       (.I0(\r_reg[2]1__2_n_65 ),
        .I1(r_reg[23]),
        .O(\n_reg[3]0_i_28__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_29 
       (.I0(\n_reg[2]0__2_n_96 ),
        .I1(\n_reg[2]0_n_96 ),
        .O(\n_reg[3]0_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_29__0 
       (.I0(\n_reg[3]0_i_48_n_7 ),
        .O(\n_reg[3]0_i_29__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_29__1 
       (.I0(\r_reg[2]1__2_n_66 ),
        .I1(r_reg[22]),
        .O(\n_reg[3]0_i_29__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_2__0 
       (.CI(\n_reg[3]0_i_3__0_n_0 ),
        .CO({\n_reg[3]0_i_2__0_n_0 ,\n_reg[3]0_i_2__0_n_1 ,\n_reg[3]0_i_2__0_n_2 ,\n_reg[3]0_i_2__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[2]0__2_n_63 ,\n_reg[2]0__2_n_64 ,\n_reg[2]0__2_n_65 ,\n_reg[2]0__2_n_66 }),
        .O(\n_next[2] [28:25]),
        .S({\n_reg[3]0_i_13__0_n_0 ,\n_reg[3]0_i_14__0_n_0 ,\n_reg[3]0_i_15__0_n_0 ,\n_reg[3]0_i_16__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_2__1 
       (.CI(\n_reg[3]0_i_3__1_n_0 ),
        .CO({\n_reg[3]0_i_2__1_n_0 ,\n_reg[3]0_i_2__1_n_1 ,\n_reg[3]0_i_2__1_n_2 ,\n_reg[3]0_i_2__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\r_reg[2]0 [28:25]),
        .S({\n_reg[3]0_i_8__0_n_0 ,\n_reg[3]0_i_9__0_n_0 ,\n_reg[3]0_i_10__1_n_0 ,\n_reg[3]0_i_11__1_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_3 
       (.CI(\n_reg[3]0_i_4_n_0 ),
        .CO({\n_reg[3]0_i_3_n_0 ,\n_reg[3]0_i_3_n_1 ,\n_reg[3]0_i_3_n_2 ,\n_reg[3]0_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[2]0__2_n_83 ,\n_reg[2]0__2_n_84 ,\n_reg[2]0__2_n_85 ,\n_reg[2]0__2_n_86 }),
        .O(\n_next[2] [8:5]),
        .S({\n_reg[3]0_i_14_n_0 ,\n_reg[3]0_i_15_n_0 ,\n_reg[3]0_i_16_n_0 ,\n_reg[3]0_i_17_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_30 
       (.I0(\n_reg[2]0__2_n_97 ),
        .I1(\n_reg[2]0_n_97 ),
        .O(\n_reg[3]0_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_30__0 
       (.I0(\n_reg[3]0_i_49_n_4 ),
        .O(\n_reg[3]0_i_30__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_30__1 
       (.I0(\r_reg[2]1__2_n_67 ),
        .I1(r_reg[21]),
        .O(\n_reg[3]0_i_30__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_31 
       (.I0(\n_reg[2]0__2_n_98 ),
        .I1(\n_reg[2]0_n_98 ),
        .O(\n_reg[3]0_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_31__0 
       (.I0(\n_reg[3]0_i_49_n_5 ),
        .O(\n_reg[3]0_i_31__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_31__1 
       (.I0(\r_reg[2]1__2_n_68 ),
        .I1(r_reg[20]),
        .O(\n_reg[3]0_i_31__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_32 
       (.CI(\<const0>__0__0 ),
        .CO({\n_reg[3]0_i_32_n_0 ,\n_reg[3]0_i_32_n_1 ,\n_reg[3]0_i_32_n_2 ,\n_reg[3]0_i_32_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[2]0__2_n_103 ,\n_reg[2]0__2_n_104 ,\n_reg[2]0__2_n_105 ,\<const0>__0__0 }),
        .S({\n_reg[3]0_i_37_n_0 ,\n_reg[3]0_i_38_n_0 ,\n_reg[3]0_i_39_n_0 ,\n_reg[2]0__1_n_89 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_32__0 
       (.I0(\n_reg[3]0_i_49_n_6 ),
        .O(\n_reg[3]0_i_32__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_32__1 
       (.I0(\r_reg[2]1__2_n_69 ),
        .I1(r_reg[19]),
        .O(\n_reg[3]0_i_32__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_33 
       (.I0(\n_reg[2]0__2_n_99 ),
        .I1(\n_reg[2]0_n_99 ),
        .O(\n_reg[3]0_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_33__0 
       (.I0(\n_reg[3]0_i_49_n_7 ),
        .O(\n_reg[3]0_i_33__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_33__1 
       (.I0(\r_reg[2]1__2_n_70 ),
        .I1(r_reg[18]),
        .O(\n_reg[3]0_i_33__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_34 
       (.I0(\n_reg[2]0__2_n_100 ),
        .I1(\n_reg[2]0_n_100 ),
        .O(\n_reg[3]0_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_34__0 
       (.I0(\n_reg[3]0_i_50_n_4 ),
        .O(\n_reg[3]0_i_34__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_35 
       (.I0(\n_reg[2]0__2_n_101 ),
        .I1(\n_reg[2]0_n_101 ),
        .O(\n_reg[3]0_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_35__0 
       (.I0(\n_reg[3]0_i_50_n_5 ),
        .O(\n_reg[3]0_i_35__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_36 
       (.I0(\n_reg[2]0__2_n_102 ),
        .I1(\n_reg[2]0_n_102 ),
        .O(\n_reg[3]0_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_36__0 
       (.I0(\n_reg[3]0_i_50_n_6 ),
        .O(\n_reg[3]0_i_36__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_37 
       (.I0(\n_reg[2]0__2_n_103 ),
        .I1(\n_reg[2]0_n_103 ),
        .O(\n_reg[3]0_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_37__0 
       (.I0(\n_reg[3]0_i_9__1_n_7 ),
        .O(\n_reg[3]0_i_37__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_38 
       (.I0(\n_reg[2]0__2_n_104 ),
        .I1(\n_reg[2]0_n_104 ),
        .O(\n_reg[3]0_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_38__0 
       (.I0(\n_reg[3]0_i_50_n_7 ),
        .O(\n_reg[3]0_i_38__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_39 
       (.I0(\n_reg[2]0__2_n_105 ),
        .I1(\n_reg[2]0_n_105 ),
        .O(\n_reg[3]0_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_39__0 
       (.I0(\n_reg[3]0_i_9__1_n_4 ),
        .O(\n_reg[3]0_i_39__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_3__0 
       (.CI(\n_reg[3]0_i_4__0_n_0 ),
        .CO({\n_reg[3]0_i_3__0_n_0 ,\n_reg[3]0_i_3__0_n_1 ,\n_reg[3]0_i_3__0_n_2 ,\n_reg[3]0_i_3__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[2]0__2_n_67 ,\n_reg[2]0__2_n_68 ,\n_reg[2]0__2_n_69 ,\n_reg[2]0__2_n_70 }),
        .O(\n_next[2] [24:21]),
        .S({\n_reg[3]0_i_17__0_n_0 ,\n_reg[3]0_i_18__0_n_0 ,\n_reg[3]0_i_19__0_n_0 ,\n_reg[3]0_i_20__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_3__1 
       (.CI(\n_reg[3]0_i_4__1_n_0 ),
        .CO({\n_reg[3]0_i_3__1_n_0 ,\n_reg[3]0_i_3__1_n_1 ,\n_reg[3]0_i_3__1_n_2 ,\n_reg[3]0_i_3__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\r_reg[2]0 [24:21]),
        .S({\n_reg[3]0_i_12__1_n_0 ,\n_reg[3]0_i_13__1_n_0 ,\n_reg[3]0_i_14__1_n_0 ,\n_reg[3]0_i_15__1_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_4 
       (.CI(\n_reg[3]0_i_5_n_0 ),
        .CO({\n_reg[3]0_i_4_n_0 ,\n_reg[3]0_i_4_n_1 ,\n_reg[3]0_i_4_n_2 ,\n_reg[3]0_i_4_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[2]0__2_n_87 ,\n_reg[2]0__2_n_88 ,\n_reg[2]0__2_n_89 ,\n_reg[2]0__2_n_90 }),
        .O(\n_next[2] [4:1]),
        .S({\n_reg[3]0_i_18_n_0 ,\n_reg[3]0_i_19_n_0 ,\n_reg[3]0_i_20_n_0 ,\n_reg[3]0_i_21_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_40 
       (.I0(\n_reg[3]0_i_9__1_n_5 ),
        .O(\n_reg[3]0_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_41 
       (.I0(\n_reg[3]0_i_9__1_n_6 ),
        .O(\n_reg[3]0_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_42 
       (.CI(\n_reg[3]0_i_51_n_0 ),
        .CO({\n_reg[3]0_i_42_n_0 ,\n_reg[3]0_i_42_n_1 ,\n_reg[3]0_i_42_n_2 ,\n_reg[3]0_i_42_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\r_reg[2]1__2_n_91 ,\r_reg[2]1__2_n_92 ,\r_reg[2]1__2_n_93 ,\r_reg[2]1__2_n_94 }),
        .S({\n_reg[3]0_i_52_n_0 ,\n_reg[3]0_i_53_n_0 ,\n_reg[3]0_i_54_n_0 ,\n_reg[3]0_i_55_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_43 
       (.I0(\r_reg[2]1__2_n_87 ),
        .I1(r_reg[1]),
        .O(\n_reg[3]0_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_44 
       (.I0(\r_reg[2]1__2_n_88 ),
        .I1(r_reg[0]),
        .O(\n_reg[3]0_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_45 
       (.I0(\r_reg[2]1__2_n_89 ),
        .I1(\r_reg[2]1_n_89 ),
        .O(\n_reg[3]0_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_46 
       (.I0(\r_reg[2]1__2_n_90 ),
        .I1(\r_reg[2]1_n_90 ),
        .O(\n_reg[3]0_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_47 
       (.CI(\n_reg[3]0_i_48_n_0 ),
        .CO({\n_reg[3]0_i_47_n_0 ,\n_reg[3]0_i_47_n_1 ,\n_reg[3]0_i_47_n_2 ,\n_reg[3]0_i_47_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\r_reg[2]1__2_n_71 ,\r_reg[2]1__2_n_72 ,\r_reg[2]1__2_n_73 ,\r_reg[2]1__2_n_74 }),
        .O({\n_reg[3]0_i_47_n_4 ,\n_reg[3]0_i_47_n_5 ,\n_reg[3]0_i_47_n_6 ,\n_reg[3]0_i_47_n_7 }),
        .S({\n_reg[3]0_i_56_n_0 ,\n_reg[3]0_i_57_n_0 ,\n_reg[3]0_i_58_n_0 ,\n_reg[3]0_i_59_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_48 
       (.CI(\n_reg[3]0_i_49_n_0 ),
        .CO({\n_reg[3]0_i_48_n_0 ,\n_reg[3]0_i_48_n_1 ,\n_reg[3]0_i_48_n_2 ,\n_reg[3]0_i_48_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\r_reg[2]1__2_n_75 ,\r_reg[2]1__2_n_76 ,\r_reg[2]1__2_n_77 ,\r_reg[2]1__2_n_78 }),
        .O({\n_reg[3]0_i_48_n_4 ,\n_reg[3]0_i_48_n_5 ,\n_reg[3]0_i_48_n_6 ,\n_reg[3]0_i_48_n_7 }),
        .S({\n_reg[3]0_i_60_n_0 ,\n_reg[3]0_i_61_n_0 ,\n_reg[3]0_i_62_n_0 ,\n_reg[3]0_i_63_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_49 
       (.CI(\n_reg[3]0_i_50_n_0 ),
        .CO({\n_reg[3]0_i_49_n_0 ,\n_reg[3]0_i_49_n_1 ,\n_reg[3]0_i_49_n_2 ,\n_reg[3]0_i_49_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\r_reg[2]1__2_n_79 ,\r_reg[2]1__2_n_80 ,\r_reg[2]1__2_n_81 ,\r_reg[2]1__2_n_82 }),
        .O({\n_reg[3]0_i_49_n_4 ,\n_reg[3]0_i_49_n_5 ,\n_reg[3]0_i_49_n_6 ,\n_reg[3]0_i_49_n_7 }),
        .S({\n_reg[3]0_i_64_n_0 ,\n_reg[3]0_i_65_n_0 ,\n_reg[3]0_i_66_n_0 ,\n_reg[3]0_i_67_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_4__0 
       (.CI(\n_reg[3]0_i_1_n_0 ),
        .CO({\n_reg[3]0_i_4__0_n_0 ,\n_reg[3]0_i_4__0_n_1 ,\n_reg[3]0_i_4__0_n_2 ,\n_reg[3]0_i_4__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[2]0__2_n_71 ,\n_reg[2]0__2_n_72 ,\n_reg[2]0__2_n_73 ,\n_reg[2]0__2_n_74 }),
        .O(\n_next[2] [20:17]),
        .S({\n_reg[3]0_i_21__0_n_0 ,\n_reg[3]0_i_22__0_n_0 ,\n_reg[3]0_i_23__0_n_0 ,\n_reg[3]0_i_24__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_4__1 
       (.CI(\n_reg[3]0_i_5__1_n_0 ),
        .CO({\n_reg[3]0_i_4__1_n_0 ,\n_reg[3]0_i_4__1_n_1 ,\n_reg[3]0_i_4__1_n_2 ,\n_reg[3]0_i_4__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\r_reg[2]0 [20:17]),
        .S({\n_reg[3]0_i_16__1_n_0 ,\n_reg[3]0_i_17__1_n_0 ,\n_reg[3]0_i_18__1_n_0 ,\n_reg[3]0_i_19__1_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_5 
       (.CI(\n_reg[3]0_i_22_n_0 ),
        .CO({\n_reg[3]0_i_5_n_0 ,\n_reg[3]0_i_5_n_1 ,\n_reg[3]0_i_5_n_2 ,\n_reg[3]0_i_5_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[2]0__2_n_91 ,\n_reg[2]0__2_n_92 ,\n_reg[2]0__2_n_93 ,\n_reg[2]0__2_n_94 }),
        .O({\n_next[2] [0],\n_reg[3]0_i_5_n_5 ,\n_reg[3]0_i_5_n_6 ,\n_reg[3]0_i_5_n_7 }),
        .S({\n_reg[3]0_i_23_n_0 ,\n_reg[3]0_i_24_n_0 ,\n_reg[3]0_i_25_n_0 ,\n_reg[3]0_i_26_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_50 
       (.CI(\n_reg[3]0_i_9__1_n_0 ),
        .CO({\n_reg[3]0_i_50_n_0 ,\n_reg[3]0_i_50_n_1 ,\n_reg[3]0_i_50_n_2 ,\n_reg[3]0_i_50_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\r_reg[2]1__2_n_83 ,\r_reg[2]1__2_n_84 ,\r_reg[2]1__2_n_85 ,\r_reg[2]1__2_n_86 }),
        .O({\n_reg[3]0_i_50_n_4 ,\n_reg[3]0_i_50_n_5 ,\n_reg[3]0_i_50_n_6 ,\n_reg[3]0_i_50_n_7 }),
        .S({\n_reg[3]0_i_68_n_0 ,\n_reg[3]0_i_69_n_0 ,\n_reg[3]0_i_70_n_0 ,\n_reg[3]0_i_71_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_51 
       (.CI(\n_reg[3]0_i_72_n_0 ),
        .CO({\n_reg[3]0_i_51_n_0 ,\n_reg[3]0_i_51_n_1 ,\n_reg[3]0_i_51_n_2 ,\n_reg[3]0_i_51_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\r_reg[2]1__2_n_95 ,\r_reg[2]1__2_n_96 ,\r_reg[2]1__2_n_97 ,\r_reg[2]1__2_n_98 }),
        .S({\n_reg[3]0_i_73_n_0 ,\n_reg[3]0_i_74_n_0 ,\n_reg[3]0_i_75_n_0 ,\n_reg[3]0_i_76_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_52 
       (.I0(\r_reg[2]1__2_n_91 ),
        .I1(\r_reg[2]1_n_91 ),
        .O(\n_reg[3]0_i_52_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_53 
       (.I0(\r_reg[2]1__2_n_92 ),
        .I1(\r_reg[2]1_n_92 ),
        .O(\n_reg[3]0_i_53_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_54 
       (.I0(\r_reg[2]1__2_n_93 ),
        .I1(\r_reg[2]1_n_93 ),
        .O(\n_reg[3]0_i_54_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_55 
       (.I0(\r_reg[2]1__2_n_94 ),
        .I1(\r_reg[2]1_n_94 ),
        .O(\n_reg[3]0_i_55_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_56 
       (.I0(\r_reg[2]1__2_n_71 ),
        .I1(r_reg[17]),
        .O(\n_reg[3]0_i_56_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_57 
       (.I0(\r_reg[2]1__2_n_72 ),
        .I1(r_reg[16]),
        .O(\n_reg[3]0_i_57_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_58 
       (.I0(\r_reg[2]1__2_n_73 ),
        .I1(r_reg[15]),
        .O(\n_reg[3]0_i_58_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_59 
       (.I0(\r_reg[2]1__2_n_74 ),
        .I1(r_reg[14]),
        .O(\n_reg[3]0_i_59_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_5__0 
       (.I0(\n_reg[3]0_i_20__1_n_5 ),
        .O(\n_reg[3]0_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_5__1 
       (.CI(\n_reg[3]0_i_6__0_n_0 ),
        .CO({\n_reg[3]0_i_5__1_n_0 ,\n_reg[3]0_i_5__1_n_1 ,\n_reg[3]0_i_5__1_n_2 ,\n_reg[3]0_i_5__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\r_reg[2]0 [16:13]),
        .S({\n_reg[3]0_i_25__0_n_0 ,\n_reg[3]0_i_26__0_n_0 ,\n_reg[3]0_i_27__0_n_0 ,\n_reg[3]0_i_28__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_6 
       (.I0(\n_reg[2]0__2_n_75 ),
        .I1(\n_reg[2]0__0_n_92 ),
        .O(\n_reg[3]0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_60 
       (.I0(\r_reg[2]1__2_n_75 ),
        .I1(r_reg[13]),
        .O(\n_reg[3]0_i_60_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_61 
       (.I0(\r_reg[2]1__2_n_76 ),
        .I1(r_reg[12]),
        .O(\n_reg[3]0_i_61_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_62 
       (.I0(\r_reg[2]1__2_n_77 ),
        .I1(r_reg[11]),
        .O(\n_reg[3]0_i_62_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_63 
       (.I0(\r_reg[2]1__2_n_78 ),
        .I1(r_reg[10]),
        .O(\n_reg[3]0_i_63_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_64 
       (.I0(\r_reg[2]1__2_n_79 ),
        .I1(r_reg[9]),
        .O(\n_reg[3]0_i_64_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_65 
       (.I0(\r_reg[2]1__2_n_80 ),
        .I1(r_reg[8]),
        .O(\n_reg[3]0_i_65_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_66 
       (.I0(\r_reg[2]1__2_n_81 ),
        .I1(r_reg[7]),
        .O(\n_reg[3]0_i_66_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_67 
       (.I0(\r_reg[2]1__2_n_82 ),
        .I1(r_reg[6]),
        .O(\n_reg[3]0_i_67_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_68 
       (.I0(\r_reg[2]1__2_n_83 ),
        .I1(r_reg[5]),
        .O(\n_reg[3]0_i_68_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_69 
       (.I0(\r_reg[2]1__2_n_84 ),
        .I1(r_reg[4]),
        .O(\n_reg[3]0_i_69_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_6__0 
       (.CI(\n_reg[3]0_i_7__1_n_0 ),
        .CO({\n_reg[3]0_i_6__0_n_0 ,\n_reg[3]0_i_6__0_n_1 ,\n_reg[3]0_i_6__0_n_2 ,\n_reg[3]0_i_6__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\r_reg[2]0 [12:9]),
        .S({\n_reg[3]0_i_29__0_n_0 ,\n_reg[3]0_i_30__0_n_0 ,\n_reg[3]0_i_31__0_n_0 ,\n_reg[3]0_i_32__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_7 
       (.I0(\n_reg[2]0__2_n_76 ),
        .I1(\n_reg[2]0__0_n_93 ),
        .O(\n_reg[3]0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_70 
       (.I0(\r_reg[2]1__2_n_85 ),
        .I1(r_reg[3]),
        .O(\n_reg[3]0_i_70_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_71 
       (.I0(\r_reg[2]1__2_n_86 ),
        .I1(r_reg[2]),
        .O(\n_reg[3]0_i_71_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_72 
       (.CI(\n_reg[3]0_i_77_n_0 ),
        .CO({\n_reg[3]0_i_72_n_0 ,\n_reg[3]0_i_72_n_1 ,\n_reg[3]0_i_72_n_2 ,\n_reg[3]0_i_72_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\r_reg[2]1__2_n_99 ,\r_reg[2]1__2_n_100 ,\r_reg[2]1__2_n_101 ,\r_reg[2]1__2_n_102 }),
        .S({\n_reg[3]0_i_78_n_0 ,\n_reg[3]0_i_79_n_0 ,\n_reg[3]0_i_80_n_0 ,\n_reg[3]0_i_81_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_73 
       (.I0(\r_reg[2]1__2_n_95 ),
        .I1(\r_reg[2]1_n_95 ),
        .O(\n_reg[3]0_i_73_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_74 
       (.I0(\r_reg[2]1__2_n_96 ),
        .I1(\r_reg[2]1_n_96 ),
        .O(\n_reg[3]0_i_74_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_75 
       (.I0(\r_reg[2]1__2_n_97 ),
        .I1(\r_reg[2]1_n_97 ),
        .O(\n_reg[3]0_i_75_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_76 
       (.I0(\r_reg[2]1__2_n_98 ),
        .I1(\r_reg[2]1_n_98 ),
        .O(\n_reg[3]0_i_76_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_77 
       (.CI(\<const0>__0__0 ),
        .CO({\n_reg[3]0_i_77_n_0 ,\n_reg[3]0_i_77_n_1 ,\n_reg[3]0_i_77_n_2 ,\n_reg[3]0_i_77_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\r_reg[2]1__2_n_103 ,\r_reg[2]1__2_n_104 ,\r_reg[2]1__2_n_105 ,\<const0>__0__0 }),
        .S({\n_reg[3]0_i_82_n_0 ,\n_reg[3]0_i_83_n_0 ,\n_reg[3]0_i_84_n_0 ,\r_reg[2]1__1_n_89 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_78 
       (.I0(\r_reg[2]1__2_n_99 ),
        .I1(\r_reg[2]1_n_99 ),
        .O(\n_reg[3]0_i_78_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_79 
       (.I0(\r_reg[2]1__2_n_100 ),
        .I1(\r_reg[2]1_n_100 ),
        .O(\n_reg[3]0_i_79_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_7__0 
       (.I0(\n_reg[3]0_i_20__1_n_6 ),
        .O(\n_reg[3]0_i_7__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_7__1 
       (.CI(\n_reg[3]0_i_8__1_n_0 ),
        .CO({\n_reg[3]0_i_7__1_n_0 ,\n_reg[3]0_i_7__1_n_1 ,\n_reg[3]0_i_7__1_n_2 ,\n_reg[3]0_i_7__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\r_reg[2]0 [8:5]),
        .S({\n_reg[3]0_i_33__0_n_0 ,\n_reg[3]0_i_34__0_n_0 ,\n_reg[3]0_i_35__0_n_0 ,\n_reg[3]0_i_36__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_8 
       (.I0(\n_reg[2]0__2_n_77 ),
        .I1(\n_reg[2]0__0_n_94 ),
        .O(\n_reg[3]0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_80 
       (.I0(\r_reg[2]1__2_n_101 ),
        .I1(\r_reg[2]1_n_101 ),
        .O(\n_reg[3]0_i_80_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_81 
       (.I0(\r_reg[2]1__2_n_102 ),
        .I1(\r_reg[2]1_n_102 ),
        .O(\n_reg[3]0_i_81_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_82 
       (.I0(\r_reg[2]1__2_n_103 ),
        .I1(\r_reg[2]1_n_103 ),
        .O(\n_reg[3]0_i_82_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_83 
       (.I0(\r_reg[2]1__2_n_104 ),
        .I1(\r_reg[2]1_n_104 ),
        .O(\n_reg[3]0_i_83_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_84 
       (.I0(\r_reg[2]1__2_n_105 ),
        .I1(\r_reg[2]1_n_105 ),
        .O(\n_reg[3]0_i_84_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_8__0 
       (.I0(\n_reg[3]0_i_20__1_n_7 ),
        .O(\n_reg[3]0_i_8__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_8__1 
       (.CI(\<const0>__0__0 ),
        .CO({\n_reg[3]0_i_8__1_n_0 ,\n_reg[3]0_i_8__1_n_1 ,\n_reg[3]0_i_8__1_n_2 ,\n_reg[3]0_i_8__1_n_3 }),
        .CYINIT(\n_reg[3]0_i_37__0_n_0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\r_reg[2]0 [4:1]),
        .S({\n_reg[3]0_i_38__0_n_0 ,\n_reg[3]0_i_39__0_n_0 ,\n_reg[3]0_i_40_n_0 ,\n_reg[3]0_i_41_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \n_reg[3]0_i_9 
       (.I0(\n_reg[2]0__2_n_78 ),
        .I1(\n_reg[2]0__0_n_95 ),
        .O(\n_reg[3]0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \n_reg[3]0_i_9__0 
       (.I0(\n_reg[3]0_i_21__1_n_4 ),
        .O(\n_reg[3]0_i_9__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3]0_i_9__1 
       (.CI(\n_reg[3]0_i_42_n_0 ),
        .CO({\n_reg[3]0_i_9__1_n_0 ,\n_reg[3]0_i_9__1_n_1 ,\n_reg[3]0_i_9__1_n_2 ,\n_reg[3]0_i_9__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\r_reg[2]1__2_n_87 ,\r_reg[2]1__2_n_88 ,\r_reg[2]1__2_n_89 ,\r_reg[2]1__2_n_90 }),
        .O({\n_reg[3]0_i_9__1_n_4 ,\n_reg[3]0_i_9__1_n_5 ,\n_reg[3]0_i_9__1_n_6 ,\n_reg[3]0_i_9__1_n_7 }),
        .S({\n_reg[3]0_i_43_n_0 ,\n_reg[3]0_i_44_n_0 ,\n_reg[3]0_i_45_n_0 ,\n_reg[3]0_i_46_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [0]),
        .Q(Z[0]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3][0]_i_1 
       (.CI(\n_reg[3][0]_i_2_n_0 ),
        .CO({\n_reg[3][0]_i_1_n_0 ,\n_reg[3][0]_i_1_n_1 ,\n_reg[3][0]_i_1_n_2 ,\n_reg[3][0]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[3]0__2_n_91 ,\n_reg[3]0__2_n_92 ,\n_reg[3]0__2_n_93 ,\n_reg[3]0__2_n_94 }),
        .O({\n_next[3] [0],\n_reg[3][0]_i_1_n_5 ,\n_reg[3][0]_i_1_n_6 ,\n_reg[3][0]_i_1_n_7 }),
        .S({\n[3][0]_i_3_n_0 ,\n[3][0]_i_4_n_0 ,\n[3][0]_i_5_n_0 ,\n[3][0]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3][0]_i_12 
       (.CI(\<const0>__0__0 ),
        .CO({\n_reg[3][0]_i_12_n_0 ,\n_reg[3][0]_i_12_n_1 ,\n_reg[3][0]_i_12_n_2 ,\n_reg[3][0]_i_12_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[3]0__2_n_103 ,\n_reg[3]0__2_n_104 ,\n_reg[3]0__2_n_105 ,\<const0>__0__0 }),
        .S({\n[3][0]_i_17_n_0 ,\n[3][0]_i_18_n_0 ,\n[3][0]_i_19_n_0 ,\n_reg[3]0__1_n_89 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3][0]_i_2 
       (.CI(\n_reg[3][0]_i_7_n_0 ),
        .CO({\n_reg[3][0]_i_2_n_0 ,\n_reg[3][0]_i_2_n_1 ,\n_reg[3][0]_i_2_n_2 ,\n_reg[3][0]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[3]0__2_n_95 ,\n_reg[3]0__2_n_96 ,\n_reg[3]0__2_n_97 ,\n_reg[3]0__2_n_98 }),
        .S({\n[3][0]_i_8_n_0 ,\n[3][0]_i_9_n_0 ,n,\n[3][0]_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3][0]_i_7 
       (.CI(\n_reg[3][0]_i_12_n_0 ),
        .CO({\n_reg[3][0]_i_7_n_0 ,\n_reg[3][0]_i_7_n_1 ,\n_reg[3][0]_i_7_n_2 ,\n_reg[3][0]_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[3]0__2_n_99 ,\n_reg[3]0__2_n_100 ,\n_reg[3]0__2_n_101 ,\n_reg[3]0__2_n_102 }),
        .S({\n[3][0]_i_13_n_0 ,\n[3][0]_i_14_n_0 ,\n[3][0]_i_15_n_0 ,\n[3][0]_i_16_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [10]),
        .Q(Z[10]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [11]),
        .Q(Z[11]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [12]),
        .Q(Z[12]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3][12]_i_1 
       (.CI(\n_reg[3][8]_i_1_n_0 ),
        .CO({\n_reg[3][12]_i_1_n_0 ,\n_reg[3][12]_i_1_n_1 ,\n_reg[3][12]_i_1_n_2 ,\n_reg[3][12]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[3]0__2_n_79 ,\n_reg[3]0__2_n_80 ,\n_reg[3]0__2_n_81 ,\n_reg[3]0__2_n_82 }),
        .O(\n_next[3] [12:9]),
        .S({\n[3][12]_i_2_n_0 ,\n[3][12]_i_3_n_0 ,\n[3][12]_i_4_n_0 ,\n[3][12]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [13]),
        .Q(Z[13]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [14]),
        .Q(Z[14]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [15]),
        .Q(Z[15]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [16]),
        .Q(Z[16]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3][16]_i_1 
       (.CI(\n_reg[3][12]_i_1_n_0 ),
        .CO({\n_reg[3][16]_i_1_n_0 ,\n_reg[3][16]_i_1_n_1 ,\n_reg[3][16]_i_1_n_2 ,\n_reg[3][16]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[3]0__2_n_75 ,\n_reg[3]0__2_n_76 ,\n_reg[3]0__2_n_77 ,\n_reg[3]0__2_n_78 }),
        .O(\n_next[3] [16:13]),
        .S({\n[3][16]_i_2_n_0 ,\n[3][16]_i_3_n_0 ,\n[3][16]_i_4_n_0 ,\n[3][16]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [17]),
        .Q(Z[17]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [18]),
        .Q(Z[18]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [19]),
        .Q(Z[19]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [1]),
        .Q(Z[1]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [20]),
        .Q(Z[20]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3][20]_i_1 
       (.CI(\n_reg[3][16]_i_1_n_0 ),
        .CO({\n_reg[3][20]_i_1_n_0 ,\n_reg[3][20]_i_1_n_1 ,\n_reg[3][20]_i_1_n_2 ,\n_reg[3][20]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[3]0__2_n_71 ,\n_reg[3]0__2_n_72 ,\n_reg[3]0__2_n_73 ,\n_reg[3]0__2_n_74 }),
        .O(\n_next[3] [20:17]),
        .S({\n[3][20]_i_2_n_0 ,\n[3][20]_i_3_n_0 ,\n[3][20]_i_4_n_0 ,\n[3][20]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [21]),
        .Q(Z[21]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [22]),
        .Q(Z[22]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [23]),
        .Q(Z[23]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [24]),
        .Q(Z[24]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3][24]_i_1 
       (.CI(\n_reg[3][20]_i_1_n_0 ),
        .CO({\n_reg[3][24]_i_1_n_0 ,\n_reg[3][24]_i_1_n_1 ,\n_reg[3][24]_i_1_n_2 ,\n_reg[3][24]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[3]0__2_n_67 ,\n_reg[3]0__2_n_68 ,\n_reg[3]0__2_n_69 ,\n_reg[3]0__2_n_70 }),
        .O(\n_next[3] [24:21]),
        .S({\n[3][24]_i_2_n_0 ,\n[3][24]_i_3_n_0 ,\n[3][24]_i_4_n_0 ,\n[3][24]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [25]),
        .Q(Z[25]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [26]),
        .Q(Z[26]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [27]),
        .Q(Z[27]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [28]),
        .Q(Z[28]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3][28]_i_1 
       (.CI(\n_reg[3][24]_i_1_n_0 ),
        .CO({\n_reg[3][28]_i_1_n_0 ,\n_reg[3][28]_i_1_n_1 ,\n_reg[3][28]_i_1_n_2 ,\n_reg[3][28]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[3]0__2_n_63 ,\n_reg[3]0__2_n_64 ,\n_reg[3]0__2_n_65 ,\n_reg[3]0__2_n_66 }),
        .O(\n_next[3] [28:25]),
        .S({\n[3][28]_i_2_n_0 ,\n[3][28]_i_3_n_0 ,\n[3][28]_i_4_n_0 ,\n[3][28]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [29]),
        .Q(Z[29]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [2]),
        .Q(Z[2]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [30]),
        .Q(Z[30]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [31]),
        .Q(Z[31]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3][31]_i_2 
       (.CI(\n_reg[3][28]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\n_reg[3]0__2_n_61 ,\n_reg[3]0__2_n_62 }),
        .O({\n_reg[3][31]_i_2_n_4 ,\n_next[3] [31:29]}),
        .S({\<const0>__0__0 ,\n[3][31]_i_3_n_0 ,\n[3][31]_i_4_n_0 ,\n[3][31]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [3]),
        .Q(Z[3]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [4]),
        .Q(Z[4]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3][4]_i_1 
       (.CI(\n_reg[3][0]_i_1_n_0 ),
        .CO({\n_reg[3][4]_i_1_n_0 ,\n_reg[3][4]_i_1_n_1 ,\n_reg[3][4]_i_1_n_2 ,\n_reg[3][4]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[3]0__2_n_87 ,\n_reg[3]0__2_n_88 ,\n_reg[3]0__2_n_89 ,\n_reg[3]0__2_n_90 }),
        .O(\n_next[3] [4:1]),
        .S({\n[3][4]_i_2_n_0 ,\n[3][4]_i_3_n_0 ,\n[3][4]_i_4_n_0 ,\n[3][4]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [5]),
        .Q(Z[5]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [6]),
        .Q(Z[6]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [7]),
        .Q(Z[7]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [8]),
        .Q(Z[8]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \n_reg[3][8]_i_1 
       (.CI(\n_reg[3][4]_i_1_n_0 ),
        .CO({\n_reg[3][8]_i_1_n_0 ,\n_reg[3][8]_i_1_n_1 ,\n_reg[3][8]_i_1_n_2 ,\n_reg[3][8]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\n_reg[3]0__2_n_83 ,\n_reg[3]0__2_n_84 ,\n_reg[3]0__2_n_85 ,\n_reg[3]0__2_n_86 }),
        .O(\n_next[3] [8:5]),
        .S({\n[3][8]_i_2_n_0 ,\n[3][8]_i_3_n_0 ,\n[3][8]_i_4_n_0 ,\n[3][8]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \n_reg[3][9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\n_next[3] [9]),
        .Q(Z[9]),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [31]),
        .Q(psdsp_n),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_1
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [30]),
        .Q(psdsp_n_1),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_10
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [21]),
        .Q(psdsp_n_10),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_11
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [20]),
        .Q(psdsp_n_11),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_12
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [19]),
        .Q(psdsp_n_12),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_13
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [18]),
        .Q(psdsp_n_13),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_14
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [17]),
        .Q(psdsp_n_14),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_15
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [31]),
        .Q(psdsp_n_15),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_16
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [30]),
        .Q(psdsp_n_16),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_17
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [29]),
        .Q(psdsp_n_17),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_18
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [28]),
        .Q(psdsp_n_18),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_19
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [27]),
        .Q(psdsp_n_19),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_2
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [29]),
        .Q(psdsp_n_2),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_20
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [26]),
        .Q(psdsp_n_20),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_21
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [25]),
        .Q(psdsp_n_21),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_22
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [24]),
        .Q(psdsp_n_22),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_23
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [23]),
        .Q(psdsp_n_23),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_24
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [22]),
        .Q(psdsp_n_24),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_25
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [21]),
        .Q(psdsp_n_25),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_26
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [20]),
        .Q(psdsp_n_26),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_27
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [19]),
        .Q(psdsp_n_27),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_28
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [18]),
        .Q(psdsp_n_28),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_29
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [17]),
        .Q(psdsp_n_29),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_3
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [28]),
        .Q(psdsp_n_3),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_30
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [16]),
        .Q(psdsp_n_30),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_31
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [15]),
        .Q(psdsp_n_31),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_32
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [14]),
        .Q(psdsp_n_32),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_33
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [13]),
        .Q(psdsp_n_33),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_34
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [12]),
        .Q(psdsp_n_34),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_35
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [11]),
        .Q(psdsp_n_35),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_36
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [10]),
        .Q(psdsp_n_36),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_37
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [9]),
        .Q(psdsp_n_37),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_38
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [8]),
        .Q(psdsp_n_38),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_39
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [7]),
        .Q(psdsp_n_39),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_4
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [27]),
        .Q(psdsp_n_4),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_40
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [6]),
        .Q(psdsp_n_40),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_41
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [5]),
        .Q(psdsp_n_41),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_42
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [4]),
        .Q(psdsp_n_42),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_43
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [3]),
        .Q(psdsp_n_43),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_44
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [2]),
        .Q(psdsp_n_44),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_45
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [1]),
        .Q(psdsp_n_45),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_46
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [0]),
        .Q(psdsp_n_46),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_47
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [16]),
        .Q(psdsp_n_47),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_48
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [15]),
        .Q(psdsp_n_48),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_49
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [14]),
        .Q(psdsp_n_49),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_5
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [26]),
        .Q(psdsp_n_5),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_50
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [13]),
        .Q(psdsp_n_50),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_51
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [12]),
        .Q(psdsp_n_51),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_52
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [11]),
        .Q(psdsp_n_52),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_53
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [10]),
        .Q(psdsp_n_53),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_54
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [9]),
        .Q(psdsp_n_54),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_55
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [8]),
        .Q(psdsp_n_55),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_56
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [7]),
        .Q(psdsp_n_56),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_57
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [6]),
        .Q(psdsp_n_57),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_58
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [5]),
        .Q(psdsp_n_58),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_59
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [4]),
        .Q(psdsp_n_59),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_6
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [25]),
        .Q(psdsp_n_6),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_60
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [3]),
        .Q(psdsp_n_60),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_61
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [2]),
        .Q(psdsp_n_61),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_62
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [1]),
        .Q(psdsp_n_62),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_63
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [0]),
        .Q(psdsp_n_63),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_7
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [24]),
        .Q(psdsp_n_7),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_8
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [23]),
        .Q(psdsp_n_8),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    psdsp_9
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\rsqr_next[1] [22]),
        .Q(psdsp_n_9),
        .R(RSTA));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-10 {cell *THIS*} {string 16x18 4}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(1),
    .BREG(1),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \r_reg[2]1 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,psdsp_n_30,psdsp_n_31,psdsp_n_32,psdsp_n_33,psdsp_n_34,psdsp_n_35,psdsp_n_36,psdsp_n_37,psdsp_n_38,psdsp_n_39,psdsp_n_40,psdsp_n_41,psdsp_n_42,psdsp_n_43,psdsp_n_44,psdsp_n_45,psdsp_n_46}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\d_next[1] [31:17]}),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const1>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const1>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\r_reg[2]1_n_58 ,\r_reg[2]1_n_59 ,\r_reg[2]1_n_60 ,\r_reg[2]1_n_61 ,\r_reg[2]1_n_62 ,\r_reg[2]1_n_63 ,\r_reg[2]1_n_64 ,\r_reg[2]1_n_65 ,\r_reg[2]1_n_66 ,\r_reg[2]1_n_67 ,\r_reg[2]1_n_68 ,\r_reg[2]1_n_69 ,\r_reg[2]1_n_70 ,\r_reg[2]1_n_71 ,\r_reg[2]1_n_72 ,\r_reg[2]1_n_73 ,\r_reg[2]1_n_74 ,\r_reg[2]1_n_75 ,\r_reg[2]1_n_76 ,\r_reg[2]1_n_77 ,\r_reg[2]1_n_78 ,\r_reg[2]1_n_79 ,\r_reg[2]1_n_80 ,\r_reg[2]1_n_81 ,\r_reg[2]1_n_82 ,\r_reg[2]1_n_83 ,\r_reg[2]1_n_84 ,\r_reg[2]1_n_85 ,\r_reg[2]1_n_86 ,\r_reg[2]1_n_87 ,\r_reg[2]1_n_88 ,\r_reg[2]1_n_89 ,\r_reg[2]1_n_90 ,\r_reg[2]1_n_91 ,\r_reg[2]1_n_92 ,\r_reg[2]1_n_93 ,\r_reg[2]1_n_94 ,\r_reg[2]1_n_95 ,\r_reg[2]1_n_96 ,\r_reg[2]1_n_97 ,\r_reg[2]1_n_98 ,\r_reg[2]1_n_99 ,\r_reg[2]1_n_100 ,\r_reg[2]1_n_101 ,\r_reg[2]1_n_102 ,\r_reg[2]1_n_103 ,\r_reg[2]1_n_104 ,\r_reg[2]1_n_105 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .PCOUT({\r_reg[2]1_n_106 ,\r_reg[2]1_n_107 ,\r_reg[2]1_n_108 ,\r_reg[2]1_n_109 ,\r_reg[2]1_n_110 ,\r_reg[2]1_n_111 ,\r_reg[2]1_n_112 ,\r_reg[2]1_n_113 ,\r_reg[2]1_n_114 ,\r_reg[2]1_n_115 ,\r_reg[2]1_n_116 ,\r_reg[2]1_n_117 ,\r_reg[2]1_n_118 ,\r_reg[2]1_n_119 ,\r_reg[2]1_n_120 ,\r_reg[2]1_n_121 ,\r_reg[2]1_n_122 ,\r_reg[2]1_n_123 ,\r_reg[2]1_n_124 ,\r_reg[2]1_n_125 ,\r_reg[2]1_n_126 ,\r_reg[2]1_n_127 ,\r_reg[2]1_n_128 ,\r_reg[2]1_n_129 ,\r_reg[2]1_n_130 ,\r_reg[2]1_n_131 ,\r_reg[2]1_n_132 ,\r_reg[2]1_n_133 ,\r_reg[2]1_n_134 ,\r_reg[2]1_n_135 ,\r_reg[2]1_n_136 ,\r_reg[2]1_n_137 ,\r_reg[2]1_n_138 ,\r_reg[2]1_n_139 ,\r_reg[2]1_n_140 ,\r_reg[2]1_n_141 ,\r_reg[2]1_n_142 ,\r_reg[2]1_n_143 ,\r_reg[2]1_n_144 ,\r_reg[2]1_n_145 ,\r_reg[2]1_n_146 ,\r_reg[2]1_n_147 ,\r_reg[2]1_n_148 ,\r_reg[2]1_n_149 ,\r_reg[2]1_n_150 ,\r_reg[2]1_n_151 ,\r_reg[2]1_n_152 ,\r_reg[2]1_n_153 }),
        .RSTA(RSTA),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(RSTA),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-10 {cell *THIS*} {string 16x16 4}}" *) 
  DSP48E1 #(
    .ACASCREG(1),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(1),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \r_reg[2]1__0 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\d_next[1] [31:17]}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,psdsp_n,psdsp_n_1,psdsp_n_2,psdsp_n_3,psdsp_n_4,psdsp_n_5,psdsp_n_6,psdsp_n_7,psdsp_n_8,psdsp_n_9,psdsp_n_10,psdsp_n_11,psdsp_n_12,psdsp_n_13,psdsp_n_14}),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const1>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const1>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P(r_reg),
        .PCIN({\r_reg[2]1_n_106 ,\r_reg[2]1_n_107 ,\r_reg[2]1_n_108 ,\r_reg[2]1_n_109 ,\r_reg[2]1_n_110 ,\r_reg[2]1_n_111 ,\r_reg[2]1_n_112 ,\r_reg[2]1_n_113 ,\r_reg[2]1_n_114 ,\r_reg[2]1_n_115 ,\r_reg[2]1_n_116 ,\r_reg[2]1_n_117 ,\r_reg[2]1_n_118 ,\r_reg[2]1_n_119 ,\r_reg[2]1_n_120 ,\r_reg[2]1_n_121 ,\r_reg[2]1_n_122 ,\r_reg[2]1_n_123 ,\r_reg[2]1_n_124 ,\r_reg[2]1_n_125 ,\r_reg[2]1_n_126 ,\r_reg[2]1_n_127 ,\r_reg[2]1_n_128 ,\r_reg[2]1_n_129 ,\r_reg[2]1_n_130 ,\r_reg[2]1_n_131 ,\r_reg[2]1_n_132 ,\r_reg[2]1_n_133 ,\r_reg[2]1_n_134 ,\r_reg[2]1_n_135 ,\r_reg[2]1_n_136 ,\r_reg[2]1_n_137 ,\r_reg[2]1_n_138 ,\r_reg[2]1_n_139 ,\r_reg[2]1_n_140 ,\r_reg[2]1_n_141 ,\r_reg[2]1_n_142 ,\r_reg[2]1_n_143 ,\r_reg[2]1_n_144 ,\r_reg[2]1_n_145 ,\r_reg[2]1_n_146 ,\r_reg[2]1_n_147 ,\r_reg[2]1_n_148 ,\r_reg[2]1_n_149 ,\r_reg[2]1_n_150 ,\r_reg[2]1_n_151 ,\r_reg[2]1_n_152 ,\r_reg[2]1_n_153 }),
        .RSTA(RSTA),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(RSTA),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-10 {cell *THIS*} {string 18x18 4}}" *) 
  DSP48E1 #(
    .ACASCREG(1),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(1),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \r_reg[2]1__1 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\d_next[1] [16:0]}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,psdsp_n_47,psdsp_n_48,psdsp_n_49,psdsp_n_50,psdsp_n_51,psdsp_n_52,psdsp_n_53,psdsp_n_54,psdsp_n_55,psdsp_n_56,psdsp_n_57,psdsp_n_58,psdsp_n_59,psdsp_n_60,psdsp_n_61,psdsp_n_62,psdsp_n_63}),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const1>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const1>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\r_reg[2]1__1_n_58 ,\r_reg[2]1__1_n_59 ,\r_reg[2]1__1_n_60 ,\r_reg[2]1__1_n_61 ,\r_reg[2]1__1_n_62 ,\r_reg[2]1__1_n_63 ,\r_reg[2]1__1_n_64 ,\r_reg[2]1__1_n_65 ,\r_reg[2]1__1_n_66 ,\r_reg[2]1__1_n_67 ,\r_reg[2]1__1_n_68 ,\r_reg[2]1__1_n_69 ,\r_reg[2]1__1_n_70 ,\r_reg[2]1__1_n_71 ,\r_reg[2]1__1_n_72 ,\r_reg[2]1__1_n_73 ,\r_reg[2]1__1_n_74 ,\r_reg[2]1__1_n_75 ,\r_reg[2]1__1_n_76 ,\r_reg[2]1__1_n_77 ,\r_reg[2]1__1_n_78 ,\r_reg[2]1__1_n_79 ,\r_reg[2]1__1_n_80 ,\r_reg[2]1__1_n_81 ,\r_reg[2]1__1_n_82 ,\r_reg[2]1__1_n_83 ,\r_reg[2]1__1_n_84 ,\r_reg[2]1__1_n_85 ,\r_reg[2]1__1_n_86 ,\r_reg[2]1__1_n_87 ,\r_reg[2]1__1_n_88 ,\r_reg[2]1__1_n_89 ,\r_reg[2]1__1_n_90 ,\r_reg[2]1__1_n_91 ,\r_reg[2]1__1_n_92 ,\r_reg[2]1__1_n_93 ,\r_reg[2]1__1_n_94 ,\r_reg[2]1__1_n_95 ,\r_reg[2]1__1_n_96 ,\r_reg[2]1__1_n_97 ,\r_reg[2]1__1_n_98 ,\r_reg[2]1__1_n_99 ,\r_reg[2]1__1_n_100 ,\r_reg[2]1__1_n_101 ,\r_reg[2]1__1_n_102 ,\r_reg[2]1__1_n_103 ,\r_reg[2]1__1_n_104 ,\r_reg[2]1__1_n_105 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .PCOUT({\r_reg[2]1__1_n_106 ,\r_reg[2]1__1_n_107 ,\r_reg[2]1__1_n_108 ,\r_reg[2]1__1_n_109 ,\r_reg[2]1__1_n_110 ,\r_reg[2]1__1_n_111 ,\r_reg[2]1__1_n_112 ,\r_reg[2]1__1_n_113 ,\r_reg[2]1__1_n_114 ,\r_reg[2]1__1_n_115 ,\r_reg[2]1__1_n_116 ,\r_reg[2]1__1_n_117 ,\r_reg[2]1__1_n_118 ,\r_reg[2]1__1_n_119 ,\r_reg[2]1__1_n_120 ,\r_reg[2]1__1_n_121 ,\r_reg[2]1__1_n_122 ,\r_reg[2]1__1_n_123 ,\r_reg[2]1__1_n_124 ,\r_reg[2]1__1_n_125 ,\r_reg[2]1__1_n_126 ,\r_reg[2]1__1_n_127 ,\r_reg[2]1__1_n_128 ,\r_reg[2]1__1_n_129 ,\r_reg[2]1__1_n_130 ,\r_reg[2]1__1_n_131 ,\r_reg[2]1__1_n_132 ,\r_reg[2]1__1_n_133 ,\r_reg[2]1__1_n_134 ,\r_reg[2]1__1_n_135 ,\r_reg[2]1__1_n_136 ,\r_reg[2]1__1_n_137 ,\r_reg[2]1__1_n_138 ,\r_reg[2]1__1_n_139 ,\r_reg[2]1__1_n_140 ,\r_reg[2]1__1_n_141 ,\r_reg[2]1__1_n_142 ,\r_reg[2]1__1_n_143 ,\r_reg[2]1__1_n_144 ,\r_reg[2]1__1_n_145 ,\r_reg[2]1__1_n_146 ,\r_reg[2]1__1_n_147 ,\r_reg[2]1__1_n_148 ,\r_reg[2]1__1_n_149 ,\r_reg[2]1__1_n_150 ,\r_reg[2]1__1_n_151 ,\r_reg[2]1__1_n_152 ,\r_reg[2]1__1_n_153 }),
        .RSTA(RSTA),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(RSTA),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-10 {cell *THIS*} {string 18x16 4}}" *) 
  DSP48E1 #(
    .ACASCREG(1),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(1),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \r_reg[2]1__2 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\d_next[1] [16:0]}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,psdsp_n_15,psdsp_n_16,psdsp_n_17,psdsp_n_18,psdsp_n_19,psdsp_n_20,psdsp_n_21,psdsp_n_22,psdsp_n_23,psdsp_n_24,psdsp_n_25,psdsp_n_26,psdsp_n_27,psdsp_n_28,psdsp_n_29}),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const1>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const1>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\r_reg[2]1__2_n_58 ,\r_reg[2]1__2_n_59 ,\r_reg[2]1__2_n_60 ,\r_reg[2]1__2_n_61 ,\r_reg[2]1__2_n_62 ,\r_reg[2]1__2_n_63 ,\r_reg[2]1__2_n_64 ,\r_reg[2]1__2_n_65 ,\r_reg[2]1__2_n_66 ,\r_reg[2]1__2_n_67 ,\r_reg[2]1__2_n_68 ,\r_reg[2]1__2_n_69 ,\r_reg[2]1__2_n_70 ,\r_reg[2]1__2_n_71 ,\r_reg[2]1__2_n_72 ,\r_reg[2]1__2_n_73 ,\r_reg[2]1__2_n_74 ,\r_reg[2]1__2_n_75 ,\r_reg[2]1__2_n_76 ,\r_reg[2]1__2_n_77 ,\r_reg[2]1__2_n_78 ,\r_reg[2]1__2_n_79 ,\r_reg[2]1__2_n_80 ,\r_reg[2]1__2_n_81 ,\r_reg[2]1__2_n_82 ,\r_reg[2]1__2_n_83 ,\r_reg[2]1__2_n_84 ,\r_reg[2]1__2_n_85 ,\r_reg[2]1__2_n_86 ,\r_reg[2]1__2_n_87 ,\r_reg[2]1__2_n_88 ,\r_reg[2]1__2_n_89 ,\r_reg[2]1__2_n_90 ,\r_reg[2]1__2_n_91 ,\r_reg[2]1__2_n_92 ,\r_reg[2]1__2_n_93 ,\r_reg[2]1__2_n_94 ,\r_reg[2]1__2_n_95 ,\r_reg[2]1__2_n_96 ,\r_reg[2]1__2_n_97 ,\r_reg[2]1__2_n_98 ,\r_reg[2]1__2_n_99 ,\r_reg[2]1__2_n_100 ,\r_reg[2]1__2_n_101 ,\r_reg[2]1__2_n_102 ,\r_reg[2]1__2_n_103 ,\r_reg[2]1__2_n_104 ,\r_reg[2]1__2_n_105 }),
        .PCIN({\r_reg[2]1__1_n_106 ,\r_reg[2]1__1_n_107 ,\r_reg[2]1__1_n_108 ,\r_reg[2]1__1_n_109 ,\r_reg[2]1__1_n_110 ,\r_reg[2]1__1_n_111 ,\r_reg[2]1__1_n_112 ,\r_reg[2]1__1_n_113 ,\r_reg[2]1__1_n_114 ,\r_reg[2]1__1_n_115 ,\r_reg[2]1__1_n_116 ,\r_reg[2]1__1_n_117 ,\r_reg[2]1__1_n_118 ,\r_reg[2]1__1_n_119 ,\r_reg[2]1__1_n_120 ,\r_reg[2]1__1_n_121 ,\r_reg[2]1__1_n_122 ,\r_reg[2]1__1_n_123 ,\r_reg[2]1__1_n_124 ,\r_reg[2]1__1_n_125 ,\r_reg[2]1__1_n_126 ,\r_reg[2]1__1_n_127 ,\r_reg[2]1__1_n_128 ,\r_reg[2]1__1_n_129 ,\r_reg[2]1__1_n_130 ,\r_reg[2]1__1_n_131 ,\r_reg[2]1__1_n_132 ,\r_reg[2]1__1_n_133 ,\r_reg[2]1__1_n_134 ,\r_reg[2]1__1_n_135 ,\r_reg[2]1__1_n_136 ,\r_reg[2]1__1_n_137 ,\r_reg[2]1__1_n_138 ,\r_reg[2]1__1_n_139 ,\r_reg[2]1__1_n_140 ,\r_reg[2]1__1_n_141 ,\r_reg[2]1__1_n_142 ,\r_reg[2]1__1_n_143 ,\r_reg[2]1__1_n_144 ,\r_reg[2]1__1_n_145 ,\r_reg[2]1__1_n_146 ,\r_reg[2]1__1_n_147 ,\r_reg[2]1__1_n_148 ,\r_reg[2]1__1_n_149 ,\r_reg[2]1__1_n_150 ,\r_reg[2]1__1_n_151 ,\r_reg[2]1__1_n_152 ,\r_reg[2]1__1_n_153 }),
        .RSTA(RSTA),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(RSTA),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[2]1_i_1 
       (.CI(\r_reg[2]1_i_2_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\rsqr_reg[1]0__2_n_61 ,\rsqr_reg[1]0__2_n_62 }),
        .O({\r_reg[2]1_i_1_n_4 ,\rsqr_next[1] [31:29]}),
        .S({\<const0>__0__0 ,\r_reg[2]1_i_5__0_n_0 ,\r_reg[2]1_i_6__0_n_0 ,\r_reg[2]1_i_7__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_10 
       (.I0(\rsqr_reg[1]0__2_n_65 ),
        .I1(rsqr_reg[23]),
        .O(\r_reg[2]1_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_10__0 
       (.I0(p_1_in[42]),
        .I1(d_reg[8]),
        .O(\r_reg[2]1_i_10__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_10__1 
       (.I0(p_1_in[62]),
        .I1(d_reg[28]),
        .O(\r_reg[2]1_i_10__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_11 
       (.I0(\rsqr_reg[1]0__2_n_66 ),
        .I1(rsqr_reg[22]),
        .O(\r_reg[2]1_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_11__0 
       (.I0(p_1_in[41]),
        .I1(d_reg[7]),
        .O(\r_reg[2]1_i_11__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_11__1 
       (.I0(p_1_in[61]),
        .I1(d_reg[27]),
        .O(\r_reg[2]1_i_11__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_12 
       (.I0(\rsqr_reg[1]0__2_n_67 ),
        .I1(rsqr_reg[21]),
        .O(\r_reg[2]1_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_12__0 
       (.I0(p_1_in[40]),
        .I1(d_reg[6]),
        .O(\r_reg[2]1_i_12__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_12__1 
       (.I0(p_1_in[60]),
        .I1(d_reg[26]),
        .O(\r_reg[2]1_i_12__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_13 
       (.I0(\rsqr_reg[1]0__2_n_68 ),
        .I1(rsqr_reg[20]),
        .O(\r_reg[2]1_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_13__0 
       (.I0(p_1_in[39]),
        .I1(d_reg[5]),
        .O(\r_reg[2]1_i_13__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_13__1 
       (.I0(p_1_in[59]),
        .I1(d_reg[25]),
        .O(\r_reg[2]1_i_13__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_14 
       (.I0(\rsqr_reg[1]0__2_n_69 ),
        .I1(rsqr_reg[19]),
        .O(\r_reg[2]1_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_14__0 
       (.I0(p_1_in[38]),
        .I1(d_reg[4]),
        .O(\r_reg[2]1_i_14__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_14__1 
       (.I0(p_1_in[58]),
        .I1(d_reg[24]),
        .O(\r_reg[2]1_i_14__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_15 
       (.I0(\rsqr_reg[1]0__2_n_70 ),
        .I1(rsqr_reg[18]),
        .O(\r_reg[2]1_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_15__0 
       (.I0(p_1_in[37]),
        .I1(d_reg[3]),
        .O(\r_reg[2]1_i_15__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_15__1 
       (.I0(p_1_in[57]),
        .I1(d_reg[23]),
        .O(\r_reg[2]1_i_15__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_16 
       (.I0(\rsqr_reg[1]0__2_n_71 ),
        .I1(rsqr_reg[17]),
        .O(\r_reg[2]1_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_16__0 
       (.I0(p_1_in[36]),
        .I1(d_reg[2]),
        .O(\r_reg[2]1_i_16__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_16__1 
       (.I0(p_1_in[56]),
        .I1(d_reg[22]),
        .O(\r_reg[2]1_i_16__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_17 
       (.I0(\rsqr_reg[1]0__2_n_72 ),
        .I1(rsqr_reg[16]),
        .O(\r_reg[2]1_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[2]1_i_17__0 
       (.CI(\r_reg[2]1_i_22_n_0 ),
        .CO({\r_reg[2]1_i_17__0_n_0 ,\r_reg[2]1_i_17__0_n_1 ,\r_reg[2]1_i_17__0_n_2 ,\r_reg[2]1_i_17__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(p_1_in[27:24]),
        .S({\r_reg[2]1_i_23_n_0 ,\r_reg[2]1_i_24_n_0 ,\r_reg[2]1_i_25__0_n_0 ,\r_reg[2]1_i_26__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_17__1 
       (.I0(p_1_in[55]),
        .I1(d_reg[21]),
        .O(\r_reg[2]1_i_17__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_18 
       (.I0(\rsqr_reg[1]0__2_n_73 ),
        .I1(rsqr_reg[15]),
        .O(\r_reg[2]1_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_18__0 
       (.I0(p_1_in[31]),
        .I1(\d_reg[1]0_n_91 ),
        .O(\r_reg[2]1_i_18__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_18__1 
       (.I0(p_1_in[54]),
        .I1(d_reg[20]),
        .O(\r_reg[2]1_i_18__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_19 
       (.I0(\rsqr_reg[1]0__2_n_74 ),
        .I1(rsqr_reg[14]),
        .O(\r_reg[2]1_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_19__0 
       (.I0(p_1_in[30]),
        .I1(\d_reg[1]0_n_92 ),
        .O(\r_reg[2]1_i_19__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_19__1 
       (.I0(p_1_in[53]),
        .I1(d_reg[19]),
        .O(\r_reg[2]1_i_19__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[2]1_i_1__0 
       (.CI(\r_reg[2]1_i_2__0_n_0 ),
        .CO({\r_reg[2]1_i_1__0_n_0 ,\r_reg[2]1_i_1__0_n_1 ,\r_reg[2]1_i_1__0_n_2 ,\r_reg[2]1_i_1__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(p_1_in[47:44]),
        .O(\d_next[1] [16:13]),
        .S({\r_reg[2]1_i_5__1_n_0 ,\r_reg[2]1_i_6__1_n_0 ,\r_reg[2]1_i_7__1_n_0 ,\r_reg[2]1_i_8__1_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[2]1_i_1__1 
       (.CI(\r_reg[2]1_i_2__1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,p_1_in[61:60]}),
        .O({\r_reg[2]1_i_1__1_n_4 ,\d_next[1] [31:29]}),
        .S({\<const0>__0__0 ,\r_reg[2]1_i_10__1_n_0 ,\r_reg[2]1_i_11__1_n_0 ,\r_reg[2]1_i_12__1_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[2]1_i_2 
       (.CI(\r_reg[2]1_i_3_n_0 ),
        .CO({\r_reg[2]1_i_2_n_0 ,\r_reg[2]1_i_2_n_1 ,\r_reg[2]1_i_2_n_2 ,\r_reg[2]1_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\rsqr_reg[1]0__2_n_63 ,\rsqr_reg[1]0__2_n_64 ,\rsqr_reg[1]0__2_n_65 ,\rsqr_reg[1]0__2_n_66 }),
        .O(\rsqr_next[1] [28:25]),
        .S({\r_reg[2]1_i_8__0_n_0 ,\r_reg[2]1_i_9__0_n_0 ,\r_reg[2]1_i_10_n_0 ,\r_reg[2]1_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_20 
       (.I0(p_1_in[29]),
        .I1(\d_reg[1]0_n_93 ),
        .O(\r_reg[2]1_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_20__0 
       (.I0(p_1_in[52]),
        .I1(d_reg[18]),
        .O(\r_reg[2]1_i_20__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_21 
       (.I0(p_1_in[28]),
        .I1(\d_reg[1]0_n_94 ),
        .O(\r_reg[2]1_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_21__0 
       (.I0(p_1_in[51]),
        .I1(d_reg[17]),
        .O(\r_reg[2]1_i_21__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[2]1_i_22 
       (.CI(\r_reg[2]1_i_27__0_n_0 ),
        .CO({\r_reg[2]1_i_22_n_0 ,\r_reg[2]1_i_22_n_1 ,\r_reg[2]1_i_22_n_2 ,\r_reg[2]1_i_22_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(p_1_in[23:20]),
        .S({\r_reg[2]1_i_28__0_n_0 ,\r_reg[2]1_i_29__0_n_0 ,\r_reg[2]1_i_30__0_n_0 ,\r_reg[2]1_i_31__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_22__0 
       (.I0(p_1_in[50]),
        .I1(d_reg[16]),
        .O(\r_reg[2]1_i_22__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_23 
       (.I0(p_1_in[27]),
        .I1(\d_reg[1]0_n_95 ),
        .O(\r_reg[2]1_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_23__0 
       (.I0(p_1_in[49]),
        .I1(d_reg[15]),
        .O(\r_reg[2]1_i_23__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_24 
       (.I0(p_1_in[26]),
        .I1(\d_reg[1]0_n_96 ),
        .O(\r_reg[2]1_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_24__0 
       (.I0(p_1_in[48]),
        .I1(d_reg[14]),
        .O(\r_reg[2]1_i_24__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_25 
       (.I0(\rsqr_reg[1]0__2_n_75 ),
        .I1(rsqr_reg[13]),
        .O(\r_reg[2]1_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_25__0 
       (.I0(p_1_in[25]),
        .I1(\d_reg[1]0_n_97 ),
        .O(\r_reg[2]1_i_25__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_26 
       (.I0(\rsqr_reg[1]0__2_n_76 ),
        .I1(rsqr_reg[12]),
        .O(\r_reg[2]1_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_26__0 
       (.I0(p_1_in[24]),
        .I1(\d_reg[1]0_n_98 ),
        .O(\r_reg[2]1_i_26__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_27 
       (.I0(\rsqr_reg[1]0__2_n_77 ),
        .I1(rsqr_reg[11]),
        .O(\r_reg[2]1_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[2]1_i_27__0 
       (.CI(\<const0>__0__0 ),
        .CO({\r_reg[2]1_i_27__0_n_0 ,\r_reg[2]1_i_27__0_n_1 ,\r_reg[2]1_i_27__0_n_2 ,\r_reg[2]1_i_27__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({p_1_in[19:17],\<const0>__0__0 }),
        .S({\r_reg[2]1_i_32__0_n_0 ,\r_reg[2]1_i_33__0_n_0 ,\r_reg[2]1_i_34__0_n_0 ,p_1_in[16]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_28 
       (.I0(\rsqr_reg[1]0__2_n_78 ),
        .I1(rsqr_reg[10]),
        .O(\r_reg[2]1_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_28__0 
       (.I0(p_1_in[23]),
        .I1(\d_reg[1]0_n_99 ),
        .O(\r_reg[2]1_i_28__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_29 
       (.I0(\rsqr_reg[1]0__2_n_79 ),
        .I1(rsqr_reg[9]),
        .O(\r_reg[2]1_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_29__0 
       (.I0(p_1_in[22]),
        .I1(\d_reg[1]0_n_100 ),
        .O(\r_reg[2]1_i_29__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[2]1_i_2__0 
       (.CI(\r_reg[2]1_i_3__0_n_0 ),
        .CO({\r_reg[2]1_i_2__0_n_0 ,\r_reg[2]1_i_2__0_n_1 ,\r_reg[2]1_i_2__0_n_2 ,\r_reg[2]1_i_2__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(p_1_in[43:40]),
        .O(\d_next[1] [12:9]),
        .S({\r_reg[2]1_i_9__1_n_0 ,\r_reg[2]1_i_10__0_n_0 ,\r_reg[2]1_i_11__0_n_0 ,\r_reg[2]1_i_12__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[2]1_i_2__1 
       (.CI(\r_reg[2]1_i_3__1_n_0 ),
        .CO({\r_reg[2]1_i_2__1_n_0 ,\r_reg[2]1_i_2__1_n_1 ,\r_reg[2]1_i_2__1_n_2 ,\r_reg[2]1_i_2__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(p_1_in[59:56]),
        .O(\d_next[1] [28:25]),
        .S({\r_reg[2]1_i_13__1_n_0 ,\r_reg[2]1_i_14__1_n_0 ,\r_reg[2]1_i_15__1_n_0 ,\r_reg[2]1_i_16__1_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[2]1_i_3 
       (.CI(\r_reg[2]1_i_4_n_0 ),
        .CO({\r_reg[2]1_i_3_n_0 ,\r_reg[2]1_i_3_n_1 ,\r_reg[2]1_i_3_n_2 ,\r_reg[2]1_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\rsqr_reg[1]0__2_n_67 ,\rsqr_reg[1]0__2_n_68 ,\rsqr_reg[1]0__2_n_69 ,\rsqr_reg[1]0__2_n_70 }),
        .O(\rsqr_next[1] [24:21]),
        .S({\r_reg[2]1_i_12_n_0 ,\r_reg[2]1_i_13_n_0 ,\r_reg[2]1_i_14_n_0 ,\r_reg[2]1_i_15_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_30 
       (.I0(\rsqr_reg[1]0__2_n_80 ),
        .I1(rsqr_reg[8]),
        .O(\r_reg[2]1_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_30__0 
       (.I0(p_1_in[21]),
        .I1(\d_reg[1]0_n_101 ),
        .O(\r_reg[2]1_i_30__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_31 
       (.I0(\rsqr_reg[1]0__2_n_81 ),
        .I1(rsqr_reg[7]),
        .O(\r_reg[2]1_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_31__0 
       (.I0(p_1_in[20]),
        .I1(\d_reg[1]0_n_102 ),
        .O(\r_reg[2]1_i_31__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_32 
       (.I0(\rsqr_reg[1]0__2_n_82 ),
        .I1(rsqr_reg[6]),
        .O(\r_reg[2]1_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_32__0 
       (.I0(p_1_in[19]),
        .I1(\d_reg[1]0_n_103 ),
        .O(\r_reg[2]1_i_32__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_33 
       (.I0(\rsqr_reg[1]0__2_n_83 ),
        .I1(rsqr_reg[5]),
        .O(\r_reg[2]1_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_33__0 
       (.I0(p_1_in[18]),
        .I1(\d_reg[1]0_n_104 ),
        .O(\r_reg[2]1_i_33__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_34 
       (.I0(\rsqr_reg[1]0__2_n_84 ),
        .I1(rsqr_reg[4]),
        .O(\r_reg[2]1_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_34__0 
       (.I0(p_1_in[17]),
        .I1(\d_reg[1]0_n_105 ),
        .O(\r_reg[2]1_i_34__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_35 
       (.I0(\rsqr_reg[1]0__2_n_85 ),
        .I1(rsqr_reg[3]),
        .O(\r_reg[2]1_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_36 
       (.I0(\rsqr_reg[1]0__2_n_86 ),
        .I1(rsqr_reg[2]),
        .O(\r_reg[2]1_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_37 
       (.I0(\rsqr_reg[1]0__2_n_87 ),
        .I1(rsqr_reg[1]),
        .O(\r_reg[2]1_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_38 
       (.I0(\rsqr_reg[1]0__2_n_88 ),
        .I1(rsqr_reg[0]),
        .O(\r_reg[2]1_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_39 
       (.I0(\rsqr_reg[1]0__2_n_89 ),
        .I1(\rsqr_reg[1]0_n_89 ),
        .O(\r_reg[2]1_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[2]1_i_3__0 
       (.CI(\rsqr_reg[1]0_i_9_n_0 ),
        .CO({\r_reg[2]1_i_3__0_n_0 ,\r_reg[2]1_i_3__0_n_1 ,\r_reg[2]1_i_3__0_n_2 ,\r_reg[2]1_i_3__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(p_1_in[39:36]),
        .O(\d_next[1] [8:5]),
        .S({\r_reg[2]1_i_13__0_n_0 ,\r_reg[2]1_i_14__0_n_0 ,\r_reg[2]1_i_15__0_n_0 ,\r_reg[2]1_i_16__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[2]1_i_3__1 
       (.CI(\r_reg[2]1_i_4__1_n_0 ),
        .CO({\r_reg[2]1_i_3__1_n_0 ,\r_reg[2]1_i_3__1_n_1 ,\r_reg[2]1_i_3__1_n_2 ,\r_reg[2]1_i_3__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(p_1_in[55:52]),
        .O(\d_next[1] [24:21]),
        .S({\r_reg[2]1_i_17__1_n_0 ,\r_reg[2]1_i_18__1_n_0 ,\r_reg[2]1_i_19__1_n_0 ,\r_reg[2]1_i_20__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[2]1_i_4 
       (.CI(\r_reg[2]1_i_5_n_0 ),
        .CO({\r_reg[2]1_i_4_n_0 ,\r_reg[2]1_i_4_n_1 ,\r_reg[2]1_i_4_n_2 ,\r_reg[2]1_i_4_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\rsqr_reg[1]0__2_n_71 ,\rsqr_reg[1]0__2_n_72 ,\rsqr_reg[1]0__2_n_73 ,\rsqr_reg[1]0__2_n_74 }),
        .O(\rsqr_next[1] [20:17]),
        .S({\r_reg[2]1_i_16_n_0 ,\r_reg[2]1_i_17_n_0 ,\r_reg[2]1_i_18_n_0 ,\r_reg[2]1_i_19_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_40 
       (.I0(\rsqr_reg[1]0__2_n_90 ),
        .I1(\rsqr_reg[1]0_n_90 ),
        .O(\r_reg[2]1_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[2]1_i_41 
       (.CI(\r_reg[2]1_i_46_n_0 ),
        .CO({\r_reg[2]1_i_41_n_0 ,\r_reg[2]1_i_41_n_1 ,\r_reg[2]1_i_41_n_2 ,\r_reg[2]1_i_41_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\rsqr_reg[1]0__2_n_95 ,\rsqr_reg[1]0__2_n_96 ,\rsqr_reg[1]0__2_n_97 ,\rsqr_reg[1]0__2_n_98 }),
        .S({\r_reg[2]1_i_47_n_0 ,\r_reg[2]1_i_48_n_0 ,\r_reg[2]1_i_49_n_0 ,\r_reg[2]1_i_50_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_42 
       (.I0(\rsqr_reg[1]0__2_n_91 ),
        .I1(\rsqr_reg[1]0_n_91 ),
        .O(\r_reg[2]1_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_43 
       (.I0(\rsqr_reg[1]0__2_n_92 ),
        .I1(\rsqr_reg[1]0_n_92 ),
        .O(\r_reg[2]1_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_44 
       (.I0(\rsqr_reg[1]0__2_n_93 ),
        .I1(\rsqr_reg[1]0_n_93 ),
        .O(\r_reg[2]1_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_45 
       (.I0(\rsqr_reg[1]0__2_n_94 ),
        .I1(\rsqr_reg[1]0_n_94 ),
        .O(\r_reg[2]1_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[2]1_i_46 
       (.CI(\r_reg[2]1_i_51_n_0 ),
        .CO({\r_reg[2]1_i_46_n_0 ,\r_reg[2]1_i_46_n_1 ,\r_reg[2]1_i_46_n_2 ,\r_reg[2]1_i_46_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\rsqr_reg[1]0__2_n_99 ,\rsqr_reg[1]0__2_n_100 ,\rsqr_reg[1]0__2_n_101 ,\rsqr_reg[1]0__2_n_102 }),
        .S({\r_reg[2]1_i_52_n_0 ,\r_reg[2]1_i_53_n_0 ,\r_reg[2]1_i_54_n_0 ,\r_reg[2]1_i_55_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_47 
       (.I0(\rsqr_reg[1]0__2_n_95 ),
        .I1(\rsqr_reg[1]0_n_95 ),
        .O(\r_reg[2]1_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_48 
       (.I0(\rsqr_reg[1]0__2_n_96 ),
        .I1(\rsqr_reg[1]0_n_96 ),
        .O(\r_reg[2]1_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_49 
       (.I0(\rsqr_reg[1]0__2_n_97 ),
        .I1(\rsqr_reg[1]0_n_97 ),
        .O(\r_reg[2]1_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[2]1_i_4__0 
       (.CI(\r_reg[2]1_i_17__0_n_0 ),
        .CO({\r_reg[2]1_i_4__0_n_0 ,\r_reg[2]1_i_4__0_n_1 ,\r_reg[2]1_i_4__0_n_2 ,\r_reg[2]1_i_4__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(p_1_in[31:28]),
        .O({\d_next[1] [0],\r_reg[2]1_i_4__0_n_5 ,\r_reg[2]1_i_4__0_n_6 ,\r_reg[2]1_i_4__0_n_7 }),
        .S({\r_reg[2]1_i_18__0_n_0 ,\r_reg[2]1_i_19__0_n_0 ,\r_reg[2]1_i_20_n_0 ,\r_reg[2]1_i_21_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[2]1_i_4__1 
       (.CI(\r_reg[2]1_i_1__0_n_0 ),
        .CO({\r_reg[2]1_i_4__1_n_0 ,\r_reg[2]1_i_4__1_n_1 ,\r_reg[2]1_i_4__1_n_2 ,\r_reg[2]1_i_4__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(p_1_in[51:48]),
        .O(\d_next[1] [20:17]),
        .S({\r_reg[2]1_i_21__0_n_0 ,\r_reg[2]1_i_22__0_n_0 ,\r_reg[2]1_i_23__0_n_0 ,\r_reg[2]1_i_24__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[2]1_i_5 
       (.CI(\r_reg[2]1_i_6_n_0 ),
        .CO({\r_reg[2]1_i_5_n_0 ,\r_reg[2]1_i_5_n_1 ,\r_reg[2]1_i_5_n_2 ,\r_reg[2]1_i_5_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\rsqr_reg[1]0__2_n_75 ,\rsqr_reg[1]0__2_n_76 ,\rsqr_reg[1]0__2_n_77 ,\rsqr_reg[1]0__2_n_78 }),
        .O(\rsqr_next[1] [16:13]),
        .S({\r_reg[2]1_i_25_n_0 ,\r_reg[2]1_i_26_n_0 ,\r_reg[2]1_i_27_n_0 ,\r_reg[2]1_i_28_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_50 
       (.I0(\rsqr_reg[1]0__2_n_98 ),
        .I1(\rsqr_reg[1]0_n_98 ),
        .O(\r_reg[2]1_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[2]1_i_51 
       (.CI(\<const0>__0__0 ),
        .CO({\r_reg[2]1_i_51_n_0 ,\r_reg[2]1_i_51_n_1 ,\r_reg[2]1_i_51_n_2 ,\r_reg[2]1_i_51_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\rsqr_reg[1]0__2_n_103 ,\rsqr_reg[1]0__2_n_104 ,\rsqr_reg[1]0__2_n_105 ,\<const0>__0__0 }),
        .S({\r_reg[2]1_i_56_n_0 ,\r_reg[2]1_i_57_n_0 ,\r_reg[2]1_i_58_n_0 ,\rsqr_reg[1]0__1_n_89 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_52 
       (.I0(\rsqr_reg[1]0__2_n_99 ),
        .I1(\rsqr_reg[1]0_n_99 ),
        .O(\r_reg[2]1_i_52_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_53 
       (.I0(\rsqr_reg[1]0__2_n_100 ),
        .I1(\rsqr_reg[1]0_n_100 ),
        .O(\r_reg[2]1_i_53_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_54 
       (.I0(\rsqr_reg[1]0__2_n_101 ),
        .I1(\rsqr_reg[1]0_n_101 ),
        .O(\r_reg[2]1_i_54_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_55 
       (.I0(\rsqr_reg[1]0__2_n_102 ),
        .I1(\rsqr_reg[1]0_n_102 ),
        .O(\r_reg[2]1_i_55_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_56 
       (.I0(\rsqr_reg[1]0__2_n_103 ),
        .I1(\rsqr_reg[1]0_n_103 ),
        .O(\r_reg[2]1_i_56_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_57 
       (.I0(\rsqr_reg[1]0__2_n_104 ),
        .I1(\rsqr_reg[1]0_n_104 ),
        .O(\r_reg[2]1_i_57_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_58 
       (.I0(\rsqr_reg[1]0__2_n_105 ),
        .I1(\rsqr_reg[1]0_n_105 ),
        .O(\r_reg[2]1_i_58_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_5__0 
       (.I0(\rsqr_reg[1]0__2_n_60 ),
        .I1(rsqr_reg[28]),
        .O(\r_reg[2]1_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_5__1 
       (.I0(p_1_in[47]),
        .I1(d_reg[13]),
        .O(\r_reg[2]1_i_5__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[2]1_i_6 
       (.CI(\r_reg[2]1_i_7_n_0 ),
        .CO({\r_reg[2]1_i_6_n_0 ,\r_reg[2]1_i_6_n_1 ,\r_reg[2]1_i_6_n_2 ,\r_reg[2]1_i_6_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\rsqr_reg[1]0__2_n_79 ,\rsqr_reg[1]0__2_n_80 ,\rsqr_reg[1]0__2_n_81 ,\rsqr_reg[1]0__2_n_82 }),
        .O(\rsqr_next[1] [12:9]),
        .S({\r_reg[2]1_i_29_n_0 ,\r_reg[2]1_i_30_n_0 ,\r_reg[2]1_i_31_n_0 ,\r_reg[2]1_i_32_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_6__0 
       (.I0(\rsqr_reg[1]0__2_n_61 ),
        .I1(rsqr_reg[27]),
        .O(\r_reg[2]1_i_6__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_6__1 
       (.I0(p_1_in[46]),
        .I1(d_reg[12]),
        .O(\r_reg[2]1_i_6__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[2]1_i_7 
       (.CI(\r_reg[2]1_i_8_n_0 ),
        .CO({\r_reg[2]1_i_7_n_0 ,\r_reg[2]1_i_7_n_1 ,\r_reg[2]1_i_7_n_2 ,\r_reg[2]1_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\rsqr_reg[1]0__2_n_83 ,\rsqr_reg[1]0__2_n_84 ,\rsqr_reg[1]0__2_n_85 ,\rsqr_reg[1]0__2_n_86 }),
        .O(\rsqr_next[1] [8:5]),
        .S({\r_reg[2]1_i_33_n_0 ,\r_reg[2]1_i_34_n_0 ,\r_reg[2]1_i_35_n_0 ,\r_reg[2]1_i_36_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_7__0 
       (.I0(\rsqr_reg[1]0__2_n_62 ),
        .I1(rsqr_reg[26]),
        .O(\r_reg[2]1_i_7__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_7__1 
       (.I0(p_1_in[45]),
        .I1(d_reg[11]),
        .O(\r_reg[2]1_i_7__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[2]1_i_8 
       (.CI(\r_reg[2]1_i_9_n_0 ),
        .CO({\r_reg[2]1_i_8_n_0 ,\r_reg[2]1_i_8_n_1 ,\r_reg[2]1_i_8_n_2 ,\r_reg[2]1_i_8_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\rsqr_reg[1]0__2_n_87 ,\rsqr_reg[1]0__2_n_88 ,\rsqr_reg[1]0__2_n_89 ,\rsqr_reg[1]0__2_n_90 }),
        .O(\rsqr_next[1] [4:1]),
        .S({\r_reg[2]1_i_37_n_0 ,\r_reg[2]1_i_38_n_0 ,\r_reg[2]1_i_39_n_0 ,\r_reg[2]1_i_40_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_8__0 
       (.I0(\rsqr_reg[1]0__2_n_63 ),
        .I1(rsqr_reg[25]),
        .O(\r_reg[2]1_i_8__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_8__1 
       (.I0(p_1_in[44]),
        .I1(d_reg[10]),
        .O(\r_reg[2]1_i_8__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[2]1_i_9 
       (.CI(\r_reg[2]1_i_41_n_0 ),
        .CO({\r_reg[2]1_i_9_n_0 ,\r_reg[2]1_i_9_n_1 ,\r_reg[2]1_i_9_n_2 ,\r_reg[2]1_i_9_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\rsqr_reg[1]0__2_n_91 ,\rsqr_reg[1]0__2_n_92 ,\rsqr_reg[1]0__2_n_93 ,\rsqr_reg[1]0__2_n_94 }),
        .O({\rsqr_next[1] [0],\r_reg[2]1_i_9_n_5 ,\r_reg[2]1_i_9_n_6 ,\r_reg[2]1_i_9_n_7 }),
        .S({\r_reg[2]1_i_42_n_0 ,\r_reg[2]1_i_43_n_0 ,\r_reg[2]1_i_44_n_0 ,\r_reg[2]1_i_45_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_9__0 
       (.I0(\rsqr_reg[1]0__2_n_64 ),
        .I1(rsqr_reg[24]),
        .O(\r_reg[2]1_i_9__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_reg[2]1_i_9__1 
       (.I0(p_1_in[43]),
        .I1(d_reg[9]),
        .O(\r_reg[2]1_i_9__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-10 {cell *THIS*} {string 16x18 4}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \rsqr_reg[1]0 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\r_reg[1]0 [16:1],\d_next[1] [1]}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\r_reg[1]0 [31:17]}),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(\<const0>__0__0 ),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\rsqr_reg[1]0_n_58 ,\rsqr_reg[1]0_n_59 ,\rsqr_reg[1]0_n_60 ,\rsqr_reg[1]0_n_61 ,\rsqr_reg[1]0_n_62 ,\rsqr_reg[1]0_n_63 ,\rsqr_reg[1]0_n_64 ,\rsqr_reg[1]0_n_65 ,\rsqr_reg[1]0_n_66 ,\rsqr_reg[1]0_n_67 ,\rsqr_reg[1]0_n_68 ,\rsqr_reg[1]0_n_69 ,\rsqr_reg[1]0_n_70 ,\rsqr_reg[1]0_n_71 ,\rsqr_reg[1]0_n_72 ,\rsqr_reg[1]0_n_73 ,\rsqr_reg[1]0_n_74 ,\rsqr_reg[1]0_n_75 ,\rsqr_reg[1]0_n_76 ,\rsqr_reg[1]0_n_77 ,\rsqr_reg[1]0_n_78 ,\rsqr_reg[1]0_n_79 ,\rsqr_reg[1]0_n_80 ,\rsqr_reg[1]0_n_81 ,\rsqr_reg[1]0_n_82 ,\rsqr_reg[1]0_n_83 ,\rsqr_reg[1]0_n_84 ,\rsqr_reg[1]0_n_85 ,\rsqr_reg[1]0_n_86 ,\rsqr_reg[1]0_n_87 ,\rsqr_reg[1]0_n_88 ,\rsqr_reg[1]0_n_89 ,\rsqr_reg[1]0_n_90 ,\rsqr_reg[1]0_n_91 ,\rsqr_reg[1]0_n_92 ,\rsqr_reg[1]0_n_93 ,\rsqr_reg[1]0_n_94 ,\rsqr_reg[1]0_n_95 ,\rsqr_reg[1]0_n_96 ,\rsqr_reg[1]0_n_97 ,\rsqr_reg[1]0_n_98 ,\rsqr_reg[1]0_n_99 ,\rsqr_reg[1]0_n_100 ,\rsqr_reg[1]0_n_101 ,\rsqr_reg[1]0_n_102 ,\rsqr_reg[1]0_n_103 ,\rsqr_reg[1]0_n_104 ,\rsqr_reg[1]0_n_105 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .PCOUT({\rsqr_reg[1]0_n_106 ,\rsqr_reg[1]0_n_107 ,\rsqr_reg[1]0_n_108 ,\rsqr_reg[1]0_n_109 ,\rsqr_reg[1]0_n_110 ,\rsqr_reg[1]0_n_111 ,\rsqr_reg[1]0_n_112 ,\rsqr_reg[1]0_n_113 ,\rsqr_reg[1]0_n_114 ,\rsqr_reg[1]0_n_115 ,\rsqr_reg[1]0_n_116 ,\rsqr_reg[1]0_n_117 ,\rsqr_reg[1]0_n_118 ,\rsqr_reg[1]0_n_119 ,\rsqr_reg[1]0_n_120 ,\rsqr_reg[1]0_n_121 ,\rsqr_reg[1]0_n_122 ,\rsqr_reg[1]0_n_123 ,\rsqr_reg[1]0_n_124 ,\rsqr_reg[1]0_n_125 ,\rsqr_reg[1]0_n_126 ,\rsqr_reg[1]0_n_127 ,\rsqr_reg[1]0_n_128 ,\rsqr_reg[1]0_n_129 ,\rsqr_reg[1]0_n_130 ,\rsqr_reg[1]0_n_131 ,\rsqr_reg[1]0_n_132 ,\rsqr_reg[1]0_n_133 ,\rsqr_reg[1]0_n_134 ,\rsqr_reg[1]0_n_135 ,\rsqr_reg[1]0_n_136 ,\rsqr_reg[1]0_n_137 ,\rsqr_reg[1]0_n_138 ,\rsqr_reg[1]0_n_139 ,\rsqr_reg[1]0_n_140 ,\rsqr_reg[1]0_n_141 ,\rsqr_reg[1]0_n_142 ,\rsqr_reg[1]0_n_143 ,\rsqr_reg[1]0_n_144 ,\rsqr_reg[1]0_n_145 ,\rsqr_reg[1]0_n_146 ,\rsqr_reg[1]0_n_147 ,\rsqr_reg[1]0_n_148 ,\rsqr_reg[1]0_n_149 ,\rsqr_reg[1]0_n_150 ,\rsqr_reg[1]0_n_151 ,\rsqr_reg[1]0_n_152 ,\rsqr_reg[1]0_n_153 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-10 {cell *THIS*} {string 16x16 4}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \rsqr_reg[1]0__0 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\r_reg[1]0 [31:17]}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\r_reg[1]0 [31:17]}),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(\<const0>__0__0 ),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P(rsqr_reg),
        .PCIN({\rsqr_reg[1]0_n_106 ,\rsqr_reg[1]0_n_107 ,\rsqr_reg[1]0_n_108 ,\rsqr_reg[1]0_n_109 ,\rsqr_reg[1]0_n_110 ,\rsqr_reg[1]0_n_111 ,\rsqr_reg[1]0_n_112 ,\rsqr_reg[1]0_n_113 ,\rsqr_reg[1]0_n_114 ,\rsqr_reg[1]0_n_115 ,\rsqr_reg[1]0_n_116 ,\rsqr_reg[1]0_n_117 ,\rsqr_reg[1]0_n_118 ,\rsqr_reg[1]0_n_119 ,\rsqr_reg[1]0_n_120 ,\rsqr_reg[1]0_n_121 ,\rsqr_reg[1]0_n_122 ,\rsqr_reg[1]0_n_123 ,\rsqr_reg[1]0_n_124 ,\rsqr_reg[1]0_n_125 ,\rsqr_reg[1]0_n_126 ,\rsqr_reg[1]0_n_127 ,\rsqr_reg[1]0_n_128 ,\rsqr_reg[1]0_n_129 ,\rsqr_reg[1]0_n_130 ,\rsqr_reg[1]0_n_131 ,\rsqr_reg[1]0_n_132 ,\rsqr_reg[1]0_n_133 ,\rsqr_reg[1]0_n_134 ,\rsqr_reg[1]0_n_135 ,\rsqr_reg[1]0_n_136 ,\rsqr_reg[1]0_n_137 ,\rsqr_reg[1]0_n_138 ,\rsqr_reg[1]0_n_139 ,\rsqr_reg[1]0_n_140 ,\rsqr_reg[1]0_n_141 ,\rsqr_reg[1]0_n_142 ,\rsqr_reg[1]0_n_143 ,\rsqr_reg[1]0_n_144 ,\rsqr_reg[1]0_n_145 ,\rsqr_reg[1]0_n_146 ,\rsqr_reg[1]0_n_147 ,\rsqr_reg[1]0_n_148 ,\rsqr_reg[1]0_n_149 ,\rsqr_reg[1]0_n_150 ,\rsqr_reg[1]0_n_151 ,\rsqr_reg[1]0_n_152 ,\rsqr_reg[1]0_n_153 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-10 {cell *THIS*} {string 18x18 4}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \rsqr_reg[1]0__1 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\r_reg[1]0 [16:1],\d_next[1] [1]}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\r_reg[1]0 [16:1],\d_next[1] [1]}),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(\<const0>__0__0 ),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\rsqr_reg[1]0__1_n_58 ,\rsqr_reg[1]0__1_n_59 ,\rsqr_reg[1]0__1_n_60 ,\rsqr_reg[1]0__1_n_61 ,\rsqr_reg[1]0__1_n_62 ,\rsqr_reg[1]0__1_n_63 ,\rsqr_reg[1]0__1_n_64 ,\rsqr_reg[1]0__1_n_65 ,\rsqr_reg[1]0__1_n_66 ,\rsqr_reg[1]0__1_n_67 ,\rsqr_reg[1]0__1_n_68 ,\rsqr_reg[1]0__1_n_69 ,\rsqr_reg[1]0__1_n_70 ,\rsqr_reg[1]0__1_n_71 ,\rsqr_reg[1]0__1_n_72 ,\rsqr_reg[1]0__1_n_73 ,\rsqr_reg[1]0__1_n_74 ,\rsqr_reg[1]0__1_n_75 ,\rsqr_reg[1]0__1_n_76 ,\rsqr_reg[1]0__1_n_77 ,\rsqr_reg[1]0__1_n_78 ,\rsqr_reg[1]0__1_n_79 ,\rsqr_reg[1]0__1_n_80 ,\rsqr_reg[1]0__1_n_81 ,\rsqr_reg[1]0__1_n_82 ,\rsqr_reg[1]0__1_n_83 ,\rsqr_reg[1]0__1_n_84 ,\rsqr_reg[1]0__1_n_85 ,\rsqr_reg[1]0__1_n_86 ,\rsqr_reg[1]0__1_n_87 ,\rsqr_reg[1]0__1_n_88 ,\rsqr_reg[1]0__1_n_89 ,\rsqr_reg[1]0__1_n_90 ,\rsqr_reg[1]0__1_n_91 ,\rsqr_reg[1]0__1_n_92 ,\rsqr_reg[1]0__1_n_93 ,\rsqr_reg[1]0__1_n_94 ,\rsqr_reg[1]0__1_n_95 ,\rsqr_reg[1]0__1_n_96 ,\rsqr_reg[1]0__1_n_97 ,\rsqr_reg[1]0__1_n_98 ,\rsqr_reg[1]0__1_n_99 ,\rsqr_reg[1]0__1_n_100 ,\rsqr_reg[1]0__1_n_101 ,\rsqr_reg[1]0__1_n_102 ,\rsqr_reg[1]0__1_n_103 ,\rsqr_reg[1]0__1_n_104 ,\rsqr_reg[1]0__1_n_105 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .PCOUT({\rsqr_reg[1]0__1_n_106 ,\rsqr_reg[1]0__1_n_107 ,\rsqr_reg[1]0__1_n_108 ,\rsqr_reg[1]0__1_n_109 ,\rsqr_reg[1]0__1_n_110 ,\rsqr_reg[1]0__1_n_111 ,\rsqr_reg[1]0__1_n_112 ,\rsqr_reg[1]0__1_n_113 ,\rsqr_reg[1]0__1_n_114 ,\rsqr_reg[1]0__1_n_115 ,\rsqr_reg[1]0__1_n_116 ,\rsqr_reg[1]0__1_n_117 ,\rsqr_reg[1]0__1_n_118 ,\rsqr_reg[1]0__1_n_119 ,\rsqr_reg[1]0__1_n_120 ,\rsqr_reg[1]0__1_n_121 ,\rsqr_reg[1]0__1_n_122 ,\rsqr_reg[1]0__1_n_123 ,\rsqr_reg[1]0__1_n_124 ,\rsqr_reg[1]0__1_n_125 ,\rsqr_reg[1]0__1_n_126 ,\rsqr_reg[1]0__1_n_127 ,\rsqr_reg[1]0__1_n_128 ,\rsqr_reg[1]0__1_n_129 ,\rsqr_reg[1]0__1_n_130 ,\rsqr_reg[1]0__1_n_131 ,\rsqr_reg[1]0__1_n_132 ,\rsqr_reg[1]0__1_n_133 ,\rsqr_reg[1]0__1_n_134 ,\rsqr_reg[1]0__1_n_135 ,\rsqr_reg[1]0__1_n_136 ,\rsqr_reg[1]0__1_n_137 ,\rsqr_reg[1]0__1_n_138 ,\rsqr_reg[1]0__1_n_139 ,\rsqr_reg[1]0__1_n_140 ,\rsqr_reg[1]0__1_n_141 ,\rsqr_reg[1]0__1_n_142 ,\rsqr_reg[1]0__1_n_143 ,\rsqr_reg[1]0__1_n_144 ,\rsqr_reg[1]0__1_n_145 ,\rsqr_reg[1]0__1_n_146 ,\rsqr_reg[1]0__1_n_147 ,\rsqr_reg[1]0__1_n_148 ,\rsqr_reg[1]0__1_n_149 ,\rsqr_reg[1]0__1_n_150 ,\rsqr_reg[1]0__1_n_151 ,\rsqr_reg[1]0__1_n_152 ,\rsqr_reg[1]0__1_n_153 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-10 {cell *THIS*} {string 18x16 4}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \rsqr_reg[1]0__2 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\r_reg[1]0 [16:1],\d_next[1] [1]}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\r_reg[1]0 [31:17]}),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(\<const0>__0__0 ),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\rsqr_reg[1]0__2_n_58 ,\rsqr_reg[1]0__2_n_59 ,\rsqr_reg[1]0__2_n_60 ,\rsqr_reg[1]0__2_n_61 ,\rsqr_reg[1]0__2_n_62 ,\rsqr_reg[1]0__2_n_63 ,\rsqr_reg[1]0__2_n_64 ,\rsqr_reg[1]0__2_n_65 ,\rsqr_reg[1]0__2_n_66 ,\rsqr_reg[1]0__2_n_67 ,\rsqr_reg[1]0__2_n_68 ,\rsqr_reg[1]0__2_n_69 ,\rsqr_reg[1]0__2_n_70 ,\rsqr_reg[1]0__2_n_71 ,\rsqr_reg[1]0__2_n_72 ,\rsqr_reg[1]0__2_n_73 ,\rsqr_reg[1]0__2_n_74 ,\rsqr_reg[1]0__2_n_75 ,\rsqr_reg[1]0__2_n_76 ,\rsqr_reg[1]0__2_n_77 ,\rsqr_reg[1]0__2_n_78 ,\rsqr_reg[1]0__2_n_79 ,\rsqr_reg[1]0__2_n_80 ,\rsqr_reg[1]0__2_n_81 ,\rsqr_reg[1]0__2_n_82 ,\rsqr_reg[1]0__2_n_83 ,\rsqr_reg[1]0__2_n_84 ,\rsqr_reg[1]0__2_n_85 ,\rsqr_reg[1]0__2_n_86 ,\rsqr_reg[1]0__2_n_87 ,\rsqr_reg[1]0__2_n_88 ,\rsqr_reg[1]0__2_n_89 ,\rsqr_reg[1]0__2_n_90 ,\rsqr_reg[1]0__2_n_91 ,\rsqr_reg[1]0__2_n_92 ,\rsqr_reg[1]0__2_n_93 ,\rsqr_reg[1]0__2_n_94 ,\rsqr_reg[1]0__2_n_95 ,\rsqr_reg[1]0__2_n_96 ,\rsqr_reg[1]0__2_n_97 ,\rsqr_reg[1]0__2_n_98 ,\rsqr_reg[1]0__2_n_99 ,\rsqr_reg[1]0__2_n_100 ,\rsqr_reg[1]0__2_n_101 ,\rsqr_reg[1]0__2_n_102 ,\rsqr_reg[1]0__2_n_103 ,\rsqr_reg[1]0__2_n_104 ,\rsqr_reg[1]0__2_n_105 }),
        .PCIN({\rsqr_reg[1]0__1_n_106 ,\rsqr_reg[1]0__1_n_107 ,\rsqr_reg[1]0__1_n_108 ,\rsqr_reg[1]0__1_n_109 ,\rsqr_reg[1]0__1_n_110 ,\rsqr_reg[1]0__1_n_111 ,\rsqr_reg[1]0__1_n_112 ,\rsqr_reg[1]0__1_n_113 ,\rsqr_reg[1]0__1_n_114 ,\rsqr_reg[1]0__1_n_115 ,\rsqr_reg[1]0__1_n_116 ,\rsqr_reg[1]0__1_n_117 ,\rsqr_reg[1]0__1_n_118 ,\rsqr_reg[1]0__1_n_119 ,\rsqr_reg[1]0__1_n_120 ,\rsqr_reg[1]0__1_n_121 ,\rsqr_reg[1]0__1_n_122 ,\rsqr_reg[1]0__1_n_123 ,\rsqr_reg[1]0__1_n_124 ,\rsqr_reg[1]0__1_n_125 ,\rsqr_reg[1]0__1_n_126 ,\rsqr_reg[1]0__1_n_127 ,\rsqr_reg[1]0__1_n_128 ,\rsqr_reg[1]0__1_n_129 ,\rsqr_reg[1]0__1_n_130 ,\rsqr_reg[1]0__1_n_131 ,\rsqr_reg[1]0__1_n_132 ,\rsqr_reg[1]0__1_n_133 ,\rsqr_reg[1]0__1_n_134 ,\rsqr_reg[1]0__1_n_135 ,\rsqr_reg[1]0__1_n_136 ,\rsqr_reg[1]0__1_n_137 ,\rsqr_reg[1]0__1_n_138 ,\rsqr_reg[1]0__1_n_139 ,\rsqr_reg[1]0__1_n_140 ,\rsqr_reg[1]0__1_n_141 ,\rsqr_reg[1]0__1_n_142 ,\rsqr_reg[1]0__1_n_143 ,\rsqr_reg[1]0__1_n_144 ,\rsqr_reg[1]0__1_n_145 ,\rsqr_reg[1]0__1_n_146 ,\rsqr_reg[1]0__1_n_147 ,\rsqr_reg[1]0__1_n_148 ,\rsqr_reg[1]0__1_n_149 ,\rsqr_reg[1]0__1_n_150 ,\rsqr_reg[1]0__1_n_151 ,\rsqr_reg[1]0__1_n_152 ,\rsqr_reg[1]0__1_n_153 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rsqr_reg[1]0_i_1 
       (.CI(\rsqr_reg[1]0_i_2_n_0 ),
        .CO({\rsqr_reg[1]0_i_1_n_0 ,\r_reg[1]0 [31],\rsqr_reg[1]0_i_1_n_2 ,\rsqr_reg[1]0_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,p_0_in[30],\<const0>__0__0 }),
        .O({\rsqr_reg[1]0_i_1_n_4 ,\rsqr_reg[1]0_i_1_n_5 ,\r_reg[1]0 [30:29]}),
        .S({\<const0>__0__0 ,\<const1>__0__0 ,\d_next[1] [31],p_0_in[29]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_10 
       (.I0(\d_next[1] [31]),
        .O(p_0_in[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_12 
       (.I0(\d_next[1] [30]),
        .O(p_0_in[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_13 
       (.I0(\d_next[1] [29]),
        .O(p_0_in[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_14 
       (.I0(\d_next[1] [28]),
        .O(p_0_in[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_15 
       (.I0(\d_next[1] [27]),
        .O(p_0_in[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_16 
       (.I0(\d_next[1] [26]),
        .O(p_0_in[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_17 
       (.I0(\d_next[1] [25]),
        .O(p_0_in[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_18 
       (.I0(\d_next[1] [24]),
        .O(p_0_in[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_19 
       (.I0(\d_next[1] [23]),
        .O(p_0_in[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rsqr_reg[1]0_i_2 
       (.CI(\rsqr_reg[1]0_i_3_n_0 ),
        .CO({\rsqr_reg[1]0_i_2_n_0 ,\rsqr_reg[1]0_i_2_n_1 ,\rsqr_reg[1]0_i_2_n_2 ,\rsqr_reg[1]0_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\r_reg[1]0 [28:25]),
        .S(p_0_in[28:25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_20 
       (.I0(\d_next[1] [22]),
        .O(p_0_in[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_21 
       (.I0(\d_next[1] [21]),
        .O(p_0_in[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_22 
       (.I0(\d_next[1] [20]),
        .O(p_0_in[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_23 
       (.I0(\d_next[1] [19]),
        .O(p_0_in[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_24 
       (.I0(\d_next[1] [18]),
        .O(p_0_in[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_25 
       (.I0(\d_next[1] [17]),
        .O(p_0_in[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_26 
       (.I0(\d_next[1] [16]),
        .O(p_0_in[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_27 
       (.I0(\d_next[1] [15]),
        .O(p_0_in[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_28 
       (.I0(\d_next[1] [14]),
        .O(p_0_in[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_29 
       (.I0(\d_next[1] [13]),
        .O(p_0_in[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rsqr_reg[1]0_i_3 
       (.CI(\rsqr_reg[1]0_i_4_n_0 ),
        .CO({\rsqr_reg[1]0_i_3_n_0 ,\rsqr_reg[1]0_i_3_n_1 ,\rsqr_reg[1]0_i_3_n_2 ,\rsqr_reg[1]0_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\r_reg[1]0 [24:21]),
        .S(p_0_in[24:21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_30 
       (.I0(\d_next[1] [12]),
        .O(p_0_in[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_31 
       (.I0(\d_next[1] [11]),
        .O(p_0_in[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_32 
       (.I0(\d_next[1] [10]),
        .O(p_0_in[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_33 
       (.I0(\d_next[1] [9]),
        .O(p_0_in[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_34 
       (.I0(\d_next[1] [8]),
        .O(p_0_in[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_35 
       (.I0(\d_next[1] [7]),
        .O(p_0_in[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_36 
       (.I0(\d_next[1] [6]),
        .O(p_0_in[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_37 
       (.I0(\d_next[1] [1]),
        .O(p_0_in[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_38 
       (.I0(\d_next[1] [5]),
        .O(p_0_in[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_39 
       (.I0(\d_next[1] [4]),
        .O(p_0_in[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rsqr_reg[1]0_i_4 
       (.CI(\rsqr_reg[1]0_i_5_n_0 ),
        .CO({\rsqr_reg[1]0_i_4_n_0 ,\rsqr_reg[1]0_i_4_n_1 ,\rsqr_reg[1]0_i_4_n_2 ,\rsqr_reg[1]0_i_4_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\r_reg[1]0 [20:17]),
        .S(p_0_in[20:17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_40 
       (.I0(\d_next[1] [3]),
        .O(p_0_in[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \rsqr_reg[1]0_i_41 
       (.I0(\d_next[1] [2]),
        .O(p_0_in[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rsqr_reg[1]0_i_42 
       (.I0(p_1_in[35]),
        .I1(d_reg[1]),
        .O(\rsqr_reg[1]0_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rsqr_reg[1]0_i_43 
       (.I0(p_1_in[34]),
        .I1(d_reg[0]),
        .O(\rsqr_reg[1]0_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rsqr_reg[1]0_i_44 
       (.I0(p_1_in[33]),
        .I1(\d_reg[1]0_n_89 ),
        .O(\rsqr_reg[1]0_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \rsqr_reg[1]0_i_45 
       (.I0(p_1_in[32]),
        .I1(\d_reg[1]0_n_90 ),
        .O(\rsqr_reg[1]0_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rsqr_reg[1]0_i_5 
       (.CI(\rsqr_reg[1]0_i_6_n_0 ),
        .CO({\rsqr_reg[1]0_i_5_n_0 ,\rsqr_reg[1]0_i_5_n_1 ,\rsqr_reg[1]0_i_5_n_2 ,\rsqr_reg[1]0_i_5_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\r_reg[1]0 [16:13]),
        .S(p_0_in[16:13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rsqr_reg[1]0_i_6 
       (.CI(\rsqr_reg[1]0_i_7_n_0 ),
        .CO({\rsqr_reg[1]0_i_6_n_0 ,\rsqr_reg[1]0_i_6_n_1 ,\rsqr_reg[1]0_i_6_n_2 ,\rsqr_reg[1]0_i_6_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\r_reg[1]0 [12:9]),
        .S(p_0_in[12:9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rsqr_reg[1]0_i_7 
       (.CI(\rsqr_reg[1]0_i_8_n_0 ),
        .CO({\rsqr_reg[1]0_i_7_n_0 ,\rsqr_reg[1]0_i_7_n_1 ,\rsqr_reg[1]0_i_7_n_2 ,\rsqr_reg[1]0_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\r_reg[1]0 [8:5]),
        .S(p_0_in[8:5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rsqr_reg[1]0_i_8 
       (.CI(\<const0>__0__0 ),
        .CO({\rsqr_reg[1]0_i_8_n_0 ,\rsqr_reg[1]0_i_8_n_1 ,\rsqr_reg[1]0_i_8_n_2 ,\rsqr_reg[1]0_i_8_n_3 }),
        .CYINIT(p_0_in[0]),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\r_reg[1]0 [4:1]),
        .S(p_0_in[4:1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \rsqr_reg[1]0_i_9 
       (.CI(\r_reg[2]1_i_4__0_n_0 ),
        .CO({\rsqr_reg[1]0_i_9_n_0 ,\rsqr_reg[1]0_i_9_n_1 ,\rsqr_reg[1]0_i_9_n_2 ,\rsqr_reg[1]0_i_9_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(p_1_in[35:32]),
        .O(\d_next[1] [4:1]),
        .S({\rsqr_reg[1]0_i_42_n_0 ,\rsqr_reg[1]0_i_43_n_0 ,\rsqr_reg[1]0_i_44_n_0 ,\rsqr_reg[1]0_i_45_n_0 }));
endmodule
