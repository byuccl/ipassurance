module hight
   (rstn,
    clk,
    i_mk_rdy,
    i_mk,
    i_post_rdy,
    i_op,
    i_text_val,
    i_text_in,
    o_text_done,
    o_text_out,
    backdoor,
    o_rdy);
  output backdoor;
  input rstn;
  input clk;
  input i_mk_rdy;
  input [127:0]i_mk;
  input i_post_rdy;
  input i_op;
  input i_text_val;
  input [63:0]i_text_in;
  output o_text_done;
  output [63:0]o_text_out;
  output o_rdy;

  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const0>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const1>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire FSM_sequential_r_pstate;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_pstate[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_pstate[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_pstate[0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_pstate[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_pstate[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_pstate[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_pstate[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_pstate[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_pstate[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_pstate[2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_pstate[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_pstate[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_pstate[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_pstate[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_pstate[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_pstate[5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire clk;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b5__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b6__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [127:0]i_mk;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_mk_rdy;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_op;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_post_rdy;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:0]i_text_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_text_val;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire o_rdy;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire o_rdy_INST_0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire o_text_done;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:0]o_text_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]p_0_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:0]p_1_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_rnd_key_0x;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_52_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_53_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_54_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_55_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_57_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_58_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_59_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_60_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_61_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_62_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_63_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_64_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_65_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_66_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_67_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[3]_i_68_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_52_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_53_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_54_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_55_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_57_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_58_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_59_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_60_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_61_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_62_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_63_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_64_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_65_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_66_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_67_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_68_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_69_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_70_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_71_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x[7]_i_72_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]r_rnd_key_0x_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x_reg[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x_reg[3]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x_reg[3]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_0x_reg[3]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_rnd_key_1x;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[3]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[3]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[3]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[3]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[3]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[3]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[3]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[3]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[3]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[3]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[3]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[3]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[3]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[3]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[3]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[3]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[7]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[7]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[7]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[7]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[7]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[7]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[7]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[7]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[7]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[7]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[7]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[7]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x[7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]r_rnd_key_1x_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x_reg[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x_reg[3]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x_reg[3]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_1x_reg[3]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_rnd_key_2x;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_2x[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_2x[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_2x[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_2x[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_2x[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_2x[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_2x[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_2x[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_2x[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_2x[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_2x[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_2x[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_2x[6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_2x[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_2x[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_rnd_key_3x;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_3x[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_3x[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_3x[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_3x[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_3x[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_3x[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_3x[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_3x[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_3x[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_3x[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_3x[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_3x[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_3x[6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_3x[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rnd_key_3x[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_xf;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[16]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[17]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[18]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[19]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[20]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[21]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[22]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[23]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[24]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[24]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[25]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[25]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[26]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[26]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[27]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[27]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[28]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[28]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[29]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[29]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[30]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[30]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[32]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[33]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[34]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[35]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[35]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[35]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[35]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[35]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[35]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[35]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[36]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[37]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[38]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[39]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[39]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[39]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[39]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[39]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[39]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[39]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[39]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[3]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[40]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[41]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[42]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[43]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[44]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[45]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[46]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[47]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[48]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[49]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[50]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[51]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[52]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[53]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[54]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[55]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[55]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[56]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[56]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[57]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[57]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[58]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[58]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[59]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[59]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[60]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[60]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[61]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[61]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[62]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[62]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[63]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[63]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[63]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[63]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[63]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[63]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[7]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[7]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[7]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[7]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[7]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[7]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf[9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]r_xf_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf_reg[35]_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf_reg[35]_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf_reg[35]_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf_reg[35]_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf_reg[39]_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf_reg[39]_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf_reg[39]_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf_reg[39]_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf_reg[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf_reg[3]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf_reg[3]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf_reg[3]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf_reg[3]_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf_reg[3]_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf_reg[3]_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf_reg[3]_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf_reg[7]_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf_reg[7]_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf_reg[7]_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_xf_reg[7]_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rstn;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CONTROL/o_xf_sel2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CONTROL/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:0]\u_CONTROL/r_pstate ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CONTROL/r_pstate_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\u_CRYPTO_PATH/u_RF/w_rf_mv ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[0]0_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[0]0_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[0]0_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[0]0_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\u_CRYPTO_PATH/u_RF/w_rf_mv[1]12_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__21_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__21_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__21_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__21_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__43 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[1]1_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[1]1_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[1]1_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[1]1_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[2]0__21_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[2]0__21_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[2]0__21_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[2]0__21_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[2]0_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[2]0_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[2]0_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[2]0_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\u_CRYPTO_PATH/u_RF/w_rf_mv[3]15_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__21_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__21_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__21_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__21_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__43 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[3]1_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[3]1_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[3]1_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_CRYPTO_PATH/u_RF/w_rf_mv[3]1_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [32:0]\u_CRYPTO_PATH/w_wf_in_mux ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_0x ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_0x[7]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_0x[7]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_0x[7]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_0x[7]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_0x[7]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_0x[7]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_1x ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_1x[7]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_1x[7]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_1x[7]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_1x[7]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_1x[7]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/r_rnd_key_1x[7]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_KEY_SCHED/u_SKG/w_base ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/w_mk0x ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/w_mk1x ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/w_mk2x ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_KEY_SCHED/u_SKG/w_mk3x ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_rf_mv;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\w_rf_mv[0]0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\w_rf_mv[0]00_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[0]0__21_carry__0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[0]0__21_carry__0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[0]0__21_carry__0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[0]0__21_carry_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[0]0__21_carry_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[0]0__21_carry_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[0]0__21_carry_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[0]0_carry__0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[0]0_carry__0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[0]0_carry__0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[0]0_carry__0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[0]0_carry_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[0]0_carry_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[0]0_carry_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[0]0_carry_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[1]1__21_carry__0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[1]1__21_carry__0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[1]1__21_carry__0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[1]1__21_carry__0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[1]1__21_carry_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[1]1__21_carry_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[1]1__21_carry_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[1]1__21_carry_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[1]1_carry__0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[1]1_carry__0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[1]1_carry__0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[1]1_carry__0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[1]1_carry_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[1]1_carry_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[1]1_carry_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[1]1_carry_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\w_rf_mv[2]0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\w_rf_mv[2]01_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[2]0__21_carry__0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[2]0__21_carry__0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[2]0__21_carry__0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[2]0__21_carry__0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[2]0__21_carry_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[2]0__21_carry_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[2]0__21_carry_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[2]0__21_carry_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[2]0_carry__0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[2]0_carry__0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[2]0_carry__0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[2]0_carry__0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[2]0_carry_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[2]0_carry_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[2]0_carry_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[2]0_carry_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[3]1__21_carry_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[3]1__21_carry_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[3]1__21_carry_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[3]1__21_carry_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[3]1__21_carry_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[3]1__21_carry_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[3]1__21_carry_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[3]1__21_carry_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[3]1_carry__0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[3]1_carry__0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[3]1_carry__0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[3]1_carry__0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[3]1_carry_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[3]1_carry_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[3]1_carry_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \w_rf_mv[3]1_carry_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]w_rnd_idx;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]w_rnd_key;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]w_sk0x_tmp;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]w_sk1x_tmp;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]w_sk2x_tmp;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]w_sk3x_tmp;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_wf_post_pre;

  assign backdoor =  w_wf_post_pre ;

  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF2F2F2F2F2F2FFF2)) 
    \FSM_sequential_r_pstate[0]_i_1 
       (.I0(\FSM_sequential_r_pstate[0]_i_2_n_0 ),
        .I1(i_text_val),
        .I2(\FSM_sequential_r_pstate[0]_i_3_n_0 ),
        .I3(\FSM_sequential_r_pstate[0]_i_4_n_0 ),
        .I4(\u_CONTROL/r_pstate [4]),
        .I5(\u_CONTROL/r_pstate [1]),
        .O(FSM_sequential_r_pstate));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \FSM_sequential_r_pstate[0]_i_2 
       (.I0(\u_CONTROL/r_pstate [4]),
        .I1(\u_CONTROL/r_pstate [3]),
        .I2(i_mk_rdy),
        .I3(\u_CONTROL/r_pstate [5]),
        .I4(\u_CONTROL/r_pstate [2]),
        .O(\FSM_sequential_r_pstate[0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000F0001001E0)) 
    \FSM_sequential_r_pstate[0]_i_3 
       (.I0(\u_CONTROL/r_pstate [4]),
        .I1(\u_CONTROL/r_pstate [3]),
        .I2(i_mk_rdy),
        .I3(\u_CONTROL/r_pstate [0]),
        .I4(\u_CONTROL/r_pstate [5]),
        .I5(\u_CONTROL/r_pstate [2]),
        .O(\FSM_sequential_r_pstate[0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1454040404041515)) 
    \FSM_sequential_r_pstate[0]_i_4 
       (.I0(\u_CONTROL/r_pstate [3]),
        .I1(i_mk_rdy),
        .I2(\u_CONTROL/r_pstate [0]),
        .I3(i_post_rdy),
        .I4(\u_CONTROL/r_pstate [5]),
        .I5(\u_CONTROL/r_pstate [2]),
        .O(\FSM_sequential_r_pstate[0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF020202)) 
    \FSM_sequential_r_pstate[1]_i_1 
       (.I0(\FSM_sequential_r_pstate[1]_i_2_n_0 ),
        .I1(\u_CONTROL/r_pstate [3]),
        .I2(\u_CONTROL/r_pstate [4]),
        .I3(\FSM_sequential_r_pstate[1]_i_3_n_0 ),
        .I4(i_mk_rdy),
        .O(\FSM_sequential_r_pstate[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1011101190901010)) 
    \FSM_sequential_r_pstate[1]_i_2 
       (.I0(\u_CONTROL/r_pstate [5]),
        .I1(\u_CONTROL/r_pstate [2]),
        .I2(\u_CONTROL/r_pstate [0]),
        .I3(i_text_val),
        .I4(i_post_rdy),
        .I5(\u_CONTROL/r_pstate [1]),
        .O(\FSM_sequential_r_pstate[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000555655570000)) 
    \FSM_sequential_r_pstate[1]_i_3 
       (.I0(\u_CONTROL/r_pstate [5]),
        .I1(\u_CONTROL/r_pstate [4]),
        .I2(\u_CONTROL/r_pstate [2]),
        .I3(\u_CONTROL/r_pstate [3]),
        .I4(\u_CONTROL/r_pstate [0]),
        .I5(\u_CONTROL/r_pstate [1]),
        .O(\FSM_sequential_r_pstate[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF88888888888)) 
    \FSM_sequential_r_pstate[2]_i_1 
       (.I0(\FSM_sequential_r_pstate[2]_i_2_n_0 ),
        .I1(\u_CONTROL/r_pstate [0]),
        .I2(\FSM_sequential_r_pstate[2]_i_3_n_0 ),
        .I3(i_text_val),
        .I4(\FSM_sequential_r_pstate[2]_i_4_n_0 ),
        .I5(i_mk_rdy),
        .O(\FSM_sequential_r_pstate[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \FSM_sequential_r_pstate[2]_i_2 
       (.I0(\u_CONTROL/r_pstate [5]),
        .I1(\u_CONTROL/r_pstate [2]),
        .I2(\u_CONTROL/r_pstate [4]),
        .I3(\u_CONTROL/r_pstate [3]),
        .I4(i_post_rdy),
        .I5(\u_CONTROL/r_pstate [1]),
        .O(\FSM_sequential_r_pstate[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010000)) 
    \FSM_sequential_r_pstate[2]_i_3 
       (.I0(\u_CONTROL/r_pstate [0]),
        .I1(\u_CONTROL/r_pstate [5]),
        .I2(\u_CONTROL/r_pstate [4]),
        .I3(\u_CONTROL/r_pstate [3]),
        .I4(\u_CONTROL/r_pstate [1]),
        .O(\FSM_sequential_r_pstate[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1212121830303070)) 
    \FSM_sequential_r_pstate[2]_i_4 
       (.I0(\u_CONTROL/r_pstate [0]),
        .I1(\u_CONTROL/r_pstate [5]),
        .I2(\u_CONTROL/r_pstate [2]),
        .I3(\u_CONTROL/r_pstate [4]),
        .I4(\u_CONTROL/r_pstate [3]),
        .I5(\u_CONTROL/r_pstate [1]),
        .O(\FSM_sequential_r_pstate[2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0440404040404040)) 
    \FSM_sequential_r_pstate[3]_i_1 
       (.I0(\u_CONTROL/r_pstate [5]),
        .I1(i_mk_rdy),
        .I2(\u_CONTROL/r_pstate [3]),
        .I3(\u_CONTROL/r_pstate [2]),
        .I4(\u_CONTROL/r_pstate [1]),
        .I5(\u_CONTROL/r_pstate [0]),
        .O(\FSM_sequential_r_pstate[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \FSM_sequential_r_pstate[4]_i_1 
       (.I0(\FSM_sequential_r_pstate[4]_i_2_n_0 ),
        .I1(i_mk_rdy),
        .O(\FSM_sequential_r_pstate[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1450505050505050)) 
    \FSM_sequential_r_pstate[4]_i_2 
       (.I0(\u_CONTROL/r_pstate [5]),
        .I1(\u_CONTROL/r_pstate [0]),
        .I2(\u_CONTROL/r_pstate [4]),
        .I3(\u_CONTROL/r_pstate [1]),
        .I4(\u_CONTROL/r_pstate [3]),
        .I5(\u_CONTROL/r_pstate [2]),
        .O(\FSM_sequential_r_pstate[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \FSM_sequential_r_pstate[5]_i_1 
       (.I0(\FSM_sequential_r_pstate[5]_i_2_n_0 ),
        .I1(\u_CONTROL/r_pstate [5]),
        .I2(\FSM_sequential_r_pstate[5]_i_3_n_0 ),
        .I3(i_mk_rdy),
        .O(\FSM_sequential_r_pstate[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \FSM_sequential_r_pstate[5]_i_2 
       (.I0(\u_CONTROL/r_pstate [4]),
        .I1(\u_CONTROL/r_pstate [3]),
        .I2(\u_CONTROL/r_pstate [0]),
        .I3(\u_CONTROL/r_pstate [2]),
        .I4(\u_CONTROL/r_pstate [1]),
        .I5(i_post_rdy),
        .O(\FSM_sequential_r_pstate[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4000020200020202)) 
    \FSM_sequential_r_pstate[5]_i_3 
       (.I0(\u_CONTROL/r_pstate [5]),
        .I1(\u_CONTROL/r_pstate [4]),
        .I2(\u_CONTROL/r_pstate [3]),
        .I3(\u_CONTROL/r_pstate [0]),
        .I4(\u_CONTROL/r_pstate [2]),
        .I5(\u_CONTROL/r_pstate [1]),
        .O(\FSM_sequential_r_pstate[5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND
       (.G(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC
       (.P(\<const1>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h609996F9F0999090)) 
    g0_b0
       (.I0(w_rnd_idx[1]),
        .I1(i_op),
        .I2(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I3(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\u_KEY_SCHED/u_SKG/w_base [4]),
        .O(g0_b0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0090066F996F6699)) 
    g0_b0__0
       (.I0(w_rnd_idx[1]),
        .I1(i_op),
        .I2(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I3(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\u_KEY_SCHED/u_SKG/w_base [4]),
        .O(g0_b0__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF00996FF99690F69)) 
    g0_b1
       (.I0(w_rnd_idx[1]),
        .I1(i_op),
        .I2(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I3(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\u_KEY_SCHED/u_SKG/w_base [4]),
        .O(g0_b1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF60F6660F90FFF0)) 
    g0_b2
       (.I0(w_rnd_idx[1]),
        .I1(i_op),
        .I2(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I3(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\u_KEY_SCHED/u_SKG/w_base [4]),
        .O(g0_b2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6609F90F6F096909)) 
    g0_b4
       (.I0(w_rnd_idx[1]),
        .I1(i_op),
        .I2(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I3(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\u_KEY_SCHED/u_SKG/w_base [4]),
        .O(g0_b4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6009909669F6F609)) 
    g0_b4__0
       (.I0(w_rnd_idx[1]),
        .I1(i_op),
        .I2(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I3(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\u_KEY_SCHED/u_SKG/w_base [4]),
        .O(g0_b4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0F00F99F6966F066)) 
    g0_b5
       (.I0(w_rnd_idx[1]),
        .I1(i_op),
        .I2(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I3(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\u_KEY_SCHED/u_SKG/w_base [4]),
        .O(g0_b5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96006FF0F6606660)) 
    g0_b5__0
       (.I0(w_rnd_idx[1]),
        .I1(i_op),
        .I2(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I3(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\u_KEY_SCHED/u_SKG/w_base [4]),
        .O(g0_b5__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF669F9690699F6F)) 
    g0_b6
       (.I0(w_rnd_idx[1]),
        .I1(i_op),
        .I2(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I3(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\u_KEY_SCHED/u_SKG/w_base [4]),
        .O(g0_b6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF0600FF966F60F96)) 
    g0_b6__0
       (.I0(w_rnd_idx[1]),
        .I1(i_op),
        .I2(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I3(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\u_KEY_SCHED/u_SKG/w_base [4]),
        .O(g0_b6__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h11114446111A4449)) 
    g0_b6_i_1
       (.I0(\u_CONTROL/r_pstate [5]),
        .I1(\u_CONTROL/r_pstate [1]),
        .I2(\u_CONTROL/r_pstate [3]),
        .I3(\u_CONTROL/r_pstate [4]),
        .I4(\u_CONTROL/r_pstate [0]),
        .I5(\u_CONTROL/r_pstate [2]),
        .O(w_rnd_idx[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    g0_b6_i_2
       (.I0(i_op),
        .I1(w_rnd_idx[0]),
        .O(\u_KEY_SCHED/u_SKG/w_base [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    g0_b6_i_3
       (.I0(i_op),
        .I1(w_rnd_idx[2]),
        .O(\u_KEY_SCHED/u_SKG/w_base [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    g0_b6_i_4
       (.I0(i_op),
        .I1(w_rnd_idx[3]),
        .O(\u_KEY_SCHED/u_SKG/w_base [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    g0_b6_i_5
       (.I0(i_op),
        .I1(w_rnd_idx[4]),
        .O(\u_KEY_SCHED/u_SKG/w_base [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000200030000FFFC)) 
    g0_b6_i_6
       (.I0(\u_CONTROL/r_pstate [1]),
        .I1(\u_CONTROL/r_pstate [2]),
        .I2(\u_CONTROL/r_pstate [4]),
        .I3(\u_CONTROL/r_pstate [3]),
        .I4(\u_CONTROL/r_pstate [0]),
        .I5(\u_CONTROL/r_pstate [5]),
        .O(w_rnd_idx[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0007000799985550)) 
    g0_b6_i_7
       (.I0(\u_CONTROL/r_pstate [2]),
        .I1(\u_CONTROL/r_pstate [1]),
        .I2(\u_CONTROL/r_pstate [4]),
        .I3(\u_CONTROL/r_pstate [3]),
        .I4(\u_CONTROL/r_pstate [0]),
        .I5(\u_CONTROL/r_pstate [5]),
        .O(w_rnd_idx[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00F800F800075F01)) 
    g0_b6_i_8
       (.I0(\u_CONTROL/r_pstate [1]),
        .I1(\u_CONTROL/r_pstate [0]),
        .I2(\u_CONTROL/r_pstate [2]),
        .I3(\u_CONTROL/r_pstate [5]),
        .I4(\u_CONTROL/r_pstate [4]),
        .I5(\u_CONTROL/r_pstate [3]),
        .O(w_rnd_idx[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FFF8005F0004)) 
    g0_b6_i_9
       (.I0(\u_CONTROL/r_pstate [1]),
        .I1(\u_CONTROL/r_pstate [0]),
        .I2(\u_CONTROL/r_pstate [2]),
        .I3(\u_CONTROL/r_pstate [3]),
        .I4(\u_CONTROL/r_pstate [5]),
        .I5(\u_CONTROL/r_pstate [4]),
        .O(w_rnd_idx[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    o_rdy_INST_0
       (.I0(o_rdy_INST_0_i_1_n_0),
        .I1(i_mk_rdy),
        .O(o_rdy));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    o_rdy_INST_0_i_1
       (.I0(\u_CONTROL/r_pstate [2]),
        .I1(\u_CONTROL/r_pstate [5]),
        .I2(\u_CONTROL/r_pstate [4]),
        .I3(\u_CONTROL/r_pstate [3]),
        .I4(\u_CONTROL/r_pstate [0]),
        .I5(\u_CONTROL/r_pstate [1]),
        .O(o_rdy_INST_0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    o_text_done_INST_0
       (.I0(\u_CONTROL/p_0_in ),
        .I1(i_post_rdy),
        .O(o_text_done));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    o_text_done_INST_0_i_1
       (.I0(\u_CONTROL/r_pstate [1]),
        .I1(\u_CONTROL/r_pstate [2]),
        .I2(\u_CONTROL/r_pstate [4]),
        .I3(\u_CONTROL/r_pstate [3]),
        .I4(\u_CONTROL/r_pstate [5]),
        .I5(\u_CONTROL/r_pstate [0]),
        .O(\u_CONTROL/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_0x[0]_i_1 
       (.I0(w_sk3x_tmp[0]),
        .I1(i_op),
        .I2(w_sk0x_tmp[0]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(r_rnd_key_0x),
        .O(p_0_in[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[0]_i_2 
       (.I0(i_mk[0]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[96]),
        .O(r_rnd_key_0x));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_0x[1]_i_1 
       (.I0(w_sk3x_tmp[1]),
        .I1(i_op),
        .I2(w_sk0x_tmp[1]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_0x[1]_i_2_n_0 ),
        .O(p_0_in[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[1]_i_2 
       (.I0(i_mk[1]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[97]),
        .O(\r_rnd_key_0x[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_0x[2]_i_1 
       (.I0(w_sk3x_tmp[2]),
        .I1(i_op),
        .I2(w_sk0x_tmp[2]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_0x[2]_i_2_n_0 ),
        .O(p_0_in[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[2]_i_2 
       (.I0(i_mk[2]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[98]),
        .O(\r_rnd_key_0x[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_0x[3]_i_1 
       (.I0(w_sk3x_tmp[3]),
        .I1(i_op),
        .I2(w_sk0x_tmp[3]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_0x[3]_i_4_n_0 ),
        .O(p_0_in[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_13 
       (.I0(\r_rnd_key_0x[3]_i_37_n_0 ),
        .I1(\r_rnd_key_0x[3]_i_38_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[3]_i_39_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[3]_i_40_n_0 ),
        .O(\r_rnd_key_0x[3]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[3]_i_14 
       (.I0(\r_rnd_key_0x[3]_i_41_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[3]_i_42_n_0 ),
        .O(\r_rnd_key_0x[3]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[3]_i_15 
       (.I0(\r_rnd_key_0x[3]_i_43_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[3]_i_44_n_0 ),
        .O(\r_rnd_key_0x[3]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_16 
       (.I0(\r_rnd_key_0x[3]_i_45_n_0 ),
        .I1(\r_rnd_key_0x[3]_i_46_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[3]_i_47_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[3]_i_48_n_0 ),
        .O(\r_rnd_key_0x[3]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[3]_i_17 
       (.I0(\r_rnd_key_0x[3]_i_49_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[3]_i_50_n_0 ),
        .O(\r_rnd_key_0x[3]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[3]_i_18 
       (.I0(\r_rnd_key_0x[3]_i_51_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[3]_i_52_n_0 ),
        .O(\r_rnd_key_0x[3]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_19 
       (.I0(\r_rnd_key_0x[3]_i_53_n_0 ),
        .I1(\r_rnd_key_0x[3]_i_54_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[3]_i_55_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[3]_i_56_n_0 ),
        .O(\r_rnd_key_0x[3]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[3]_i_20 
       (.I0(\r_rnd_key_0x[3]_i_57_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[3]_i_58_n_0 ),
        .O(\r_rnd_key_0x[3]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[3]_i_21 
       (.I0(\r_rnd_key_0x[3]_i_59_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[3]_i_60_n_0 ),
        .O(\r_rnd_key_0x[3]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_22 
       (.I0(\r_rnd_key_0x[3]_i_61_n_0 ),
        .I1(\r_rnd_key_0x[3]_i_62_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[3]_i_63_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[3]_i_64_n_0 ),
        .O(\r_rnd_key_0x[3]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[3]_i_23 
       (.I0(\r_rnd_key_0x[3]_i_65_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[3]_i_66_n_0 ),
        .O(\r_rnd_key_0x[3]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[3]_i_24 
       (.I0(\r_rnd_key_0x[3]_i_67_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[3]_i_68_n_0 ),
        .O(\r_rnd_key_0x[3]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_25 
       (.I0(\r_rnd_key_0x[3]_i_44_n_0 ),
        .I1(\r_rnd_key_0x[3]_i_41_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[3]_i_42_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[3]_i_37_n_0 ),
        .O(\r_rnd_key_0x[3]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[3]_i_26 
       (.I0(\r_rnd_key_0x[3]_i_40_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[3]_i_43_n_0 ),
        .O(\r_rnd_key_0x[3]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[3]_i_27 
       (.I0(\r_rnd_key_0x[3]_i_38_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[3]_i_39_n_0 ),
        .O(\r_rnd_key_0x[3]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_28 
       (.I0(\r_rnd_key_0x[3]_i_52_n_0 ),
        .I1(\r_rnd_key_0x[3]_i_49_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[3]_i_50_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[3]_i_45_n_0 ),
        .O(\r_rnd_key_0x[3]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[3]_i_29 
       (.I0(\r_rnd_key_0x[3]_i_48_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[3]_i_51_n_0 ),
        .O(\r_rnd_key_0x[3]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[3]_i_30 
       (.I0(\r_rnd_key_0x[3]_i_46_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[3]_i_47_n_0 ),
        .O(\r_rnd_key_0x[3]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_31 
       (.I0(\r_rnd_key_0x[3]_i_60_n_0 ),
        .I1(\r_rnd_key_0x[3]_i_57_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[3]_i_58_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[3]_i_53_n_0 ),
        .O(\r_rnd_key_0x[3]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[3]_i_32 
       (.I0(\r_rnd_key_0x[3]_i_56_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[3]_i_59_n_0 ),
        .O(\r_rnd_key_0x[3]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[3]_i_33 
       (.I0(\r_rnd_key_0x[3]_i_54_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[3]_i_55_n_0 ),
        .O(\r_rnd_key_0x[3]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_34 
       (.I0(\r_rnd_key_0x[3]_i_68_n_0 ),
        .I1(\r_rnd_key_0x[3]_i_65_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[3]_i_66_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[3]_i_61_n_0 ),
        .O(\r_rnd_key_0x[3]_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[3]_i_35 
       (.I0(\r_rnd_key_0x[3]_i_64_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[3]_i_67_n_0 ),
        .O(\r_rnd_key_0x[3]_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[3]_i_36 
       (.I0(\r_rnd_key_0x[3]_i_62_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[3]_i_63_n_0 ),
        .O(\r_rnd_key_0x[3]_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_37 
       (.I0(i_mk[35]),
        .I1(i_mk[3]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[99]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[67]),
        .O(\r_rnd_key_0x[3]_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_38 
       (.I0(i_mk[43]),
        .I1(i_mk[11]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[107]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[75]),
        .O(\r_rnd_key_0x[3]_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_39 
       (.I0(i_mk[51]),
        .I1(i_mk[19]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[115]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[83]),
        .O(\r_rnd_key_0x[3]_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[3]_i_4 
       (.I0(i_mk[3]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[99]),
        .O(\r_rnd_key_0x[3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_40 
       (.I0(i_mk[59]),
        .I1(i_mk[27]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[123]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[91]),
        .O(\r_rnd_key_0x[3]_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_41 
       (.I0(i_mk[19]),
        .I1(i_mk[51]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[83]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[115]),
        .O(\r_rnd_key_0x[3]_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_42 
       (.I0(i_mk[27]),
        .I1(i_mk[59]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[91]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[123]),
        .O(\r_rnd_key_0x[3]_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_43 
       (.I0(i_mk[3]),
        .I1(i_mk[35]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[67]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[99]),
        .O(\r_rnd_key_0x[3]_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_44 
       (.I0(i_mk[11]),
        .I1(i_mk[43]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[75]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[107]),
        .O(\r_rnd_key_0x[3]_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_45 
       (.I0(i_mk[34]),
        .I1(i_mk[2]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[98]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[66]),
        .O(\r_rnd_key_0x[3]_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_46 
       (.I0(i_mk[42]),
        .I1(i_mk[10]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[106]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[74]),
        .O(\r_rnd_key_0x[3]_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_47 
       (.I0(i_mk[50]),
        .I1(i_mk[18]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[114]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[82]),
        .O(\r_rnd_key_0x[3]_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_48 
       (.I0(i_mk[58]),
        .I1(i_mk[26]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[122]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[90]),
        .O(\r_rnd_key_0x[3]_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_49 
       (.I0(i_mk[18]),
        .I1(i_mk[50]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[82]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[114]),
        .O(\r_rnd_key_0x[3]_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_50 
       (.I0(i_mk[26]),
        .I1(i_mk[58]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[90]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[122]),
        .O(\r_rnd_key_0x[3]_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_51 
       (.I0(i_mk[2]),
        .I1(i_mk[34]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[66]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[98]),
        .O(\r_rnd_key_0x[3]_i_51_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_52 
       (.I0(i_mk[10]),
        .I1(i_mk[42]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[74]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[106]),
        .O(\r_rnd_key_0x[3]_i_52_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_53 
       (.I0(i_mk[33]),
        .I1(i_mk[1]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[97]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[65]),
        .O(\r_rnd_key_0x[3]_i_53_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_54 
       (.I0(i_mk[41]),
        .I1(i_mk[9]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[105]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[73]),
        .O(\r_rnd_key_0x[3]_i_54_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_55 
       (.I0(i_mk[49]),
        .I1(i_mk[17]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[113]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[81]),
        .O(\r_rnd_key_0x[3]_i_55_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_56 
       (.I0(i_mk[57]),
        .I1(i_mk[25]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[121]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[89]),
        .O(\r_rnd_key_0x[3]_i_56_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_57 
       (.I0(i_mk[17]),
        .I1(i_mk[49]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[81]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[113]),
        .O(\r_rnd_key_0x[3]_i_57_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_58 
       (.I0(i_mk[25]),
        .I1(i_mk[57]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[89]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[121]),
        .O(\r_rnd_key_0x[3]_i_58_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_59 
       (.I0(i_mk[1]),
        .I1(i_mk[33]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[65]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[97]),
        .O(\r_rnd_key_0x[3]_i_59_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_60 
       (.I0(i_mk[9]),
        .I1(i_mk[41]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[73]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[105]),
        .O(\r_rnd_key_0x[3]_i_60_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_61 
       (.I0(i_mk[32]),
        .I1(i_mk[0]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[96]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[64]),
        .O(\r_rnd_key_0x[3]_i_61_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_62 
       (.I0(i_mk[40]),
        .I1(i_mk[8]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[104]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[72]),
        .O(\r_rnd_key_0x[3]_i_62_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_63 
       (.I0(i_mk[48]),
        .I1(i_mk[16]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[112]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[80]),
        .O(\r_rnd_key_0x[3]_i_63_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_64 
       (.I0(i_mk[56]),
        .I1(i_mk[24]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[120]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[88]),
        .O(\r_rnd_key_0x[3]_i_64_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_65 
       (.I0(i_mk[16]),
        .I1(i_mk[48]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[80]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[112]),
        .O(\r_rnd_key_0x[3]_i_65_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_66 
       (.I0(i_mk[24]),
        .I1(i_mk[56]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[88]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[120]),
        .O(\r_rnd_key_0x[3]_i_66_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_67 
       (.I0(i_mk[0]),
        .I1(i_mk[32]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[64]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[96]),
        .O(\r_rnd_key_0x[3]_i_67_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[3]_i_68 
       (.I0(i_mk[8]),
        .I1(i_mk[40]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[72]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[104]),
        .O(\r_rnd_key_0x[3]_i_68_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_0x[4]_i_1 
       (.I0(w_sk3x_tmp[4]),
        .I1(i_op),
        .I2(w_sk0x_tmp[4]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_0x[4]_i_2_n_0 ),
        .O(p_0_in[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[4]_i_2 
       (.I0(i_mk[4]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[100]),
        .O(\r_rnd_key_0x[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_0x[5]_i_1 
       (.I0(w_sk3x_tmp[5]),
        .I1(i_op),
        .I2(w_sk0x_tmp[5]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_0x[5]_i_2_n_0 ),
        .O(p_0_in[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[5]_i_2 
       (.I0(i_mk[5]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[101]),
        .O(\r_rnd_key_0x[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_0x[6]_i_1 
       (.I0(w_sk3x_tmp[6]),
        .I1(i_op),
        .I2(w_sk0x_tmp[6]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_0x[6]_i_2_n_0 ),
        .O(p_0_in[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[6]_i_2 
       (.I0(i_mk[6]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[102]),
        .O(\r_rnd_key_0x[6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_0x[7]_i_1 
       (.I0(w_sk3x_tmp[7]),
        .I1(i_op),
        .I2(w_sk0x_tmp[7]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_0x[7]_i_5_n_0 ),
        .O(p_0_in[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_10 
       (.I0(\r_rnd_key_0x[7]_i_27_n_0 ),
        .I1(\r_rnd_key_0x[7]_i_28_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[7]_i_29_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[7]_i_30_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/w_mk0x ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[7]_i_14 
       (.I0(\r_rnd_key_0x[7]_i_40_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_41_n_0 ),
        .O(\r_rnd_key_0x[7]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[7]_i_15 
       (.I0(\r_rnd_key_0x[7]_i_42_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_43_n_0 ),
        .O(\r_rnd_key_0x[7]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[7]_i_16 
       (.I0(\r_rnd_key_0x[7]_i_44_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_45_n_0 ),
        .O(\r_rnd_key_0x[7]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[7]_i_17 
       (.I0(\r_rnd_key_0x[7]_i_46_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_47_n_0 ),
        .O(\r_rnd_key_0x[7]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_18 
       (.I0(\r_rnd_key_0x[7]_i_48_n_0 ),
        .I1(\r_rnd_key_0x[7]_i_49_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[7]_i_50_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[7]_i_51_n_0 ),
        .O(\r_rnd_key_0x[7]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[7]_i_19 
       (.I0(\r_rnd_key_0x[7]_i_52_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_53_n_0 ),
        .O(\r_rnd_key_0x[7]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[7]_i_20 
       (.I0(\r_rnd_key_0x[7]_i_54_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_55_n_0 ),
        .O(\r_rnd_key_0x[7]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_21 
       (.I0(\r_rnd_key_0x[7]_i_56_n_0 ),
        .I1(\r_rnd_key_0x[7]_i_57_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[7]_i_58_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[7]_i_59_n_0 ),
        .O(\r_rnd_key_0x[7]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[7]_i_22 
       (.I0(\r_rnd_key_0x[7]_i_60_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_61_n_0 ),
        .O(\r_rnd_key_0x[7]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[7]_i_23 
       (.I0(\r_rnd_key_0x[7]_i_62_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_63_n_0 ),
        .O(\r_rnd_key_0x[7]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_24 
       (.I0(\r_rnd_key_0x[7]_i_64_n_0 ),
        .I1(\r_rnd_key_0x[7]_i_65_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[7]_i_66_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[7]_i_67_n_0 ),
        .O(\r_rnd_key_0x[7]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[7]_i_25 
       (.I0(\r_rnd_key_0x[7]_i_68_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_69_n_0 ),
        .O(\r_rnd_key_0x[7]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[7]_i_26 
       (.I0(\r_rnd_key_0x[7]_i_70_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_71_n_0 ),
        .O(\r_rnd_key_0x[7]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[7]_i_27 
       (.I0(\r_rnd_key_0x[7]_i_45_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_46_n_0 ),
        .O(\r_rnd_key_0x[7]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[7]_i_28 
       (.I0(\r_rnd_key_0x[7]_i_47_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_40_n_0 ),
        .O(\r_rnd_key_0x[7]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[7]_i_29 
       (.I0(\r_rnd_key_0x[7]_i_41_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_42_n_0 ),
        .O(\r_rnd_key_0x[7]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[7]_i_30 
       (.I0(\r_rnd_key_0x[7]_i_43_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_44_n_0 ),
        .O(\r_rnd_key_0x[7]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_31 
       (.I0(\r_rnd_key_0x[7]_i_55_n_0 ),
        .I1(\r_rnd_key_0x[7]_i_52_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[7]_i_53_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[7]_i_48_n_0 ),
        .O(\r_rnd_key_0x[7]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[7]_i_32 
       (.I0(\r_rnd_key_0x[7]_i_51_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_54_n_0 ),
        .O(\r_rnd_key_0x[7]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[7]_i_33 
       (.I0(\r_rnd_key_0x[7]_i_49_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_50_n_0 ),
        .O(\r_rnd_key_0x[7]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_34 
       (.I0(\r_rnd_key_0x[7]_i_63_n_0 ),
        .I1(\r_rnd_key_0x[7]_i_60_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[7]_i_61_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[7]_i_56_n_0 ),
        .O(\r_rnd_key_0x[7]_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[7]_i_35 
       (.I0(\r_rnd_key_0x[7]_i_59_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_62_n_0 ),
        .O(\r_rnd_key_0x[7]_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[7]_i_36 
       (.I0(\r_rnd_key_0x[7]_i_57_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_58_n_0 ),
        .O(\r_rnd_key_0x[7]_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_37 
       (.I0(\r_rnd_key_0x[7]_i_71_n_0 ),
        .I1(\r_rnd_key_0x[7]_i_68_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[7]_i_69_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[7]_i_64_n_0 ),
        .O(\r_rnd_key_0x[7]_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[7]_i_38 
       (.I0(\r_rnd_key_0x[7]_i_67_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_70_n_0 ),
        .O(\r_rnd_key_0x[7]_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[7]_i_39 
       (.I0(\r_rnd_key_0x[7]_i_65_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_66_n_0 ),
        .O(\r_rnd_key_0x[7]_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF444)) 
    \r_rnd_key_0x[7]_i_4 
       (.I0(\u_CONTROL/r_pstate_reg ),
        .I1(\r_xf[63]_i_4_n_0 ),
        .I2(i_text_val),
        .I3(o_rdy_INST_0_i_1_n_0),
        .O(\r_rnd_key_0x[7]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_40 
       (.I0(i_mk[7]),
        .I1(i_mk[39]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[71]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[103]),
        .O(\r_rnd_key_0x[7]_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_41 
       (.I0(i_mk[15]),
        .I1(i_mk[47]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[79]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[111]),
        .O(\r_rnd_key_0x[7]_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_42 
       (.I0(i_mk[23]),
        .I1(i_mk[55]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[87]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[119]),
        .O(\r_rnd_key_0x[7]_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_43 
       (.I0(i_mk[31]),
        .I1(i_mk[63]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[95]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[127]),
        .O(\r_rnd_key_0x[7]_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_44 
       (.I0(i_mk[39]),
        .I1(i_mk[7]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[103]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[71]),
        .O(\r_rnd_key_0x[7]_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_45 
       (.I0(i_mk[47]),
        .I1(i_mk[15]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[111]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[79]),
        .O(\r_rnd_key_0x[7]_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_46 
       (.I0(i_mk[55]),
        .I1(i_mk[23]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[119]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[87]),
        .O(\r_rnd_key_0x[7]_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_47 
       (.I0(i_mk[63]),
        .I1(i_mk[31]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[127]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[95]),
        .O(\r_rnd_key_0x[7]_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_48 
       (.I0(i_mk[38]),
        .I1(i_mk[6]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[102]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[70]),
        .O(\r_rnd_key_0x[7]_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_49 
       (.I0(i_mk[46]),
        .I1(i_mk[14]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[110]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[78]),
        .O(\r_rnd_key_0x[7]_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_0x[7]_i_5 
       (.I0(i_mk[7]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[103]),
        .O(\r_rnd_key_0x[7]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_50 
       (.I0(i_mk[54]),
        .I1(i_mk[22]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[118]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[86]),
        .O(\r_rnd_key_0x[7]_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_51 
       (.I0(i_mk[62]),
        .I1(i_mk[30]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[126]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[94]),
        .O(\r_rnd_key_0x[7]_i_51_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_52 
       (.I0(i_mk[22]),
        .I1(i_mk[54]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[86]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[118]),
        .O(\r_rnd_key_0x[7]_i_52_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_53 
       (.I0(i_mk[30]),
        .I1(i_mk[62]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[94]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[126]),
        .O(\r_rnd_key_0x[7]_i_53_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_54 
       (.I0(i_mk[6]),
        .I1(i_mk[38]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[70]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[102]),
        .O(\r_rnd_key_0x[7]_i_54_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_55 
       (.I0(i_mk[14]),
        .I1(i_mk[46]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[78]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[110]),
        .O(\r_rnd_key_0x[7]_i_55_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_56 
       (.I0(i_mk[37]),
        .I1(i_mk[5]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[101]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[69]),
        .O(\r_rnd_key_0x[7]_i_56_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_57 
       (.I0(i_mk[45]),
        .I1(i_mk[13]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[109]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[77]),
        .O(\r_rnd_key_0x[7]_i_57_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_58 
       (.I0(i_mk[53]),
        .I1(i_mk[21]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[117]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[85]),
        .O(\r_rnd_key_0x[7]_i_58_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_59 
       (.I0(i_mk[61]),
        .I1(i_mk[29]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[125]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[93]),
        .O(\r_rnd_key_0x[7]_i_59_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_6 
       (.I0(\r_rnd_key_0x[7]_i_14_n_0 ),
        .I1(\r_rnd_key_0x[7]_i_15_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[7]_i_16_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[7]_i_17_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/w_mk3x ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_60 
       (.I0(i_mk[21]),
        .I1(i_mk[53]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[85]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[117]),
        .O(\r_rnd_key_0x[7]_i_60_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_61 
       (.I0(i_mk[29]),
        .I1(i_mk[61]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[93]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[125]),
        .O(\r_rnd_key_0x[7]_i_61_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_62 
       (.I0(i_mk[5]),
        .I1(i_mk[37]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[69]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[101]),
        .O(\r_rnd_key_0x[7]_i_62_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_63 
       (.I0(i_mk[13]),
        .I1(i_mk[45]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[77]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[109]),
        .O(\r_rnd_key_0x[7]_i_63_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_64 
       (.I0(i_mk[36]),
        .I1(i_mk[4]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[100]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[68]),
        .O(\r_rnd_key_0x[7]_i_64_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_65 
       (.I0(i_mk[44]),
        .I1(i_mk[12]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[108]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[76]),
        .O(\r_rnd_key_0x[7]_i_65_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_66 
       (.I0(i_mk[52]),
        .I1(i_mk[20]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[116]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[84]),
        .O(\r_rnd_key_0x[7]_i_66_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_67 
       (.I0(i_mk[60]),
        .I1(i_mk[28]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[124]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[92]),
        .O(\r_rnd_key_0x[7]_i_67_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_68 
       (.I0(i_mk[20]),
        .I1(i_mk[52]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[84]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[116]),
        .O(\r_rnd_key_0x[7]_i_68_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_69 
       (.I0(i_mk[28]),
        .I1(i_mk[60]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[92]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[124]),
        .O(\r_rnd_key_0x[7]_i_69_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_70 
       (.I0(i_mk[4]),
        .I1(i_mk[36]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[68]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[100]),
        .O(\r_rnd_key_0x[7]_i_70_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_0x[7]_i_71 
       (.I0(i_mk[12]),
        .I1(i_mk[44]),
        .I2(\r_rnd_key_0x[7]_i_72_n_0 ),
        .I3(i_mk[76]),
        .I4(\u_KEY_SCHED/u_SKG/w_base [0]),
        .I5(i_mk[108]),
        .O(\r_rnd_key_0x[7]_i_71_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \r_rnd_key_0x[7]_i_72 
       (.I0(i_op),
        .I1(w_rnd_idx[1]),
        .O(\r_rnd_key_0x[7]_i_72_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_rnd_key_0x_reg[3]_i_2 
       (.CI(\<const0>__0__0 ),
        .CO(r_rnd_key_0x_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({g0_b6_n_0,g0_b5_n_0,g0_b4_n_0,g0_b0__0_n_0}),
        .O(w_sk3x_tmp[3:0]),
        .S({\u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_5_n_0 ,\u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_6_n_0 ,\u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_7_n_0 ,\u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_8_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_rnd_key_0x_reg[3]_i_3 
       (.CI(\<const0>__0__0 ),
        .CO({\r_rnd_key_0x_reg[3]_i_3_n_0 ,\r_rnd_key_0x_reg[3]_i_3_n_1 ,\r_rnd_key_0x_reg[3]_i_3_n_2 ,\r_rnd_key_0x_reg[3]_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({g0_b0__0_n_0,g0_b2_n_0,g0_b1_n_0,g0_b0_n_0}),
        .O(w_sk0x_tmp[3:0]),
        .S({\u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_9_n_0 ,\u_KEY_SCHED/u_SKG/r_rnd_key_0x ,\u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_11_n_0 ,\u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_12_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_rnd_key_0x_reg[7]_i_2 
       (.CI(r_rnd_key_0x_reg[3]),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,g0_b6__0_n_0,g0_b5__0_n_0,g0_b4__0_n_0}),
        .O(w_sk3x_tmp[7:4]),
        .S({\u_KEY_SCHED/u_SKG/w_mk3x ,\u_KEY_SCHED/u_SKG/r_rnd_key_0x[7]_i_7_n_0 ,\u_KEY_SCHED/u_SKG/r_rnd_key_0x[7]_i_8_n_0 ,\u_KEY_SCHED/u_SKG/r_rnd_key_0x[7]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_rnd_key_0x_reg[7]_i_3 
       (.CI(\r_rnd_key_0x_reg[3]_i_3_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,g0_b6_n_0,g0_b5_n_0,g0_b4_n_0}),
        .O(w_sk0x_tmp[7:4]),
        .S({\u_KEY_SCHED/u_SKG/w_mk0x ,\u_KEY_SCHED/u_SKG/r_rnd_key_0x[7]_i_11_n_0 ,\u_KEY_SCHED/u_SKG/r_rnd_key_0x[7]_i_12_n_0 ,\u_KEY_SCHED/u_SKG/r_rnd_key_0x[7]_i_13_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_1x[0]_i_1 
       (.I0(w_sk2x_tmp[0]),
        .I1(i_op),
        .I2(w_sk1x_tmp[0]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_1x[0]_i_2_n_0 ),
        .O(r_rnd_key_1x));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_1x[0]_i_2 
       (.I0(i_mk[8]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[104]),
        .O(\r_rnd_key_1x[0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_1x[1]_i_1 
       (.I0(w_sk2x_tmp[1]),
        .I1(i_op),
        .I2(w_sk1x_tmp[1]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_1x[1]_i_2_n_0 ),
        .O(\r_rnd_key_1x[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_1x[1]_i_2 
       (.I0(i_mk[9]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[105]),
        .O(\r_rnd_key_1x[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_1x[2]_i_1 
       (.I0(w_sk2x_tmp[2]),
        .I1(i_op),
        .I2(w_sk1x_tmp[2]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_1x[2]_i_2_n_0 ),
        .O(\r_rnd_key_1x[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_1x[2]_i_2 
       (.I0(i_mk[10]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[106]),
        .O(\r_rnd_key_1x[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_1x[3]_i_1 
       (.I0(w_sk2x_tmp[3]),
        .I1(i_op),
        .I2(w_sk1x_tmp[3]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_1x[3]_i_4_n_0 ),
        .O(\r_rnd_key_1x[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_1x[3]_i_13 
       (.I0(\r_rnd_key_0x[3]_i_42_n_0 ),
        .I1(\r_rnd_key_0x[3]_i_37_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[3]_i_38_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[3]_i_39_n_0 ),
        .O(\r_rnd_key_1x[3]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_1x[3]_i_14 
       (.I0(\r_rnd_key_0x[3]_i_44_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[3]_i_41_n_0 ),
        .O(\r_rnd_key_1x[3]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_1x[3]_i_15 
       (.I0(\r_rnd_key_0x[3]_i_50_n_0 ),
        .I1(\r_rnd_key_0x[3]_i_45_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[3]_i_46_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[3]_i_47_n_0 ),
        .O(\r_rnd_key_1x[3]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_1x[3]_i_16 
       (.I0(\r_rnd_key_0x[3]_i_52_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[3]_i_49_n_0 ),
        .O(\r_rnd_key_1x[3]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_1x[3]_i_17 
       (.I0(\r_rnd_key_0x[3]_i_58_n_0 ),
        .I1(\r_rnd_key_0x[3]_i_53_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[3]_i_54_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[3]_i_55_n_0 ),
        .O(\r_rnd_key_1x[3]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_1x[3]_i_18 
       (.I0(\r_rnd_key_0x[3]_i_60_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[3]_i_57_n_0 ),
        .O(\r_rnd_key_1x[3]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_1x[3]_i_19 
       (.I0(\r_rnd_key_0x[3]_i_66_n_0 ),
        .I1(\r_rnd_key_0x[3]_i_61_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[3]_i_62_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[3]_i_63_n_0 ),
        .O(\r_rnd_key_1x[3]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_1x[3]_i_20 
       (.I0(\r_rnd_key_0x[3]_i_68_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[3]_i_65_n_0 ),
        .O(\r_rnd_key_1x[3]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_1x[3]_i_21 
       (.I0(\r_rnd_key_0x[3]_i_41_n_0 ),
        .I1(\r_rnd_key_0x[3]_i_42_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[3]_i_37_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[3]_i_38_n_0 ),
        .O(\r_rnd_key_1x[3]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_1x[3]_i_22 
       (.I0(\r_rnd_key_0x[3]_i_39_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[3]_i_40_n_0 ),
        .O(\r_rnd_key_1x[3]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_1x[3]_i_23 
       (.I0(\r_rnd_key_0x[3]_i_49_n_0 ),
        .I1(\r_rnd_key_0x[3]_i_50_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[3]_i_45_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[3]_i_46_n_0 ),
        .O(\r_rnd_key_1x[3]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_1x[3]_i_24 
       (.I0(\r_rnd_key_0x[3]_i_47_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[3]_i_48_n_0 ),
        .O(\r_rnd_key_1x[3]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_1x[3]_i_25 
       (.I0(\r_rnd_key_0x[3]_i_57_n_0 ),
        .I1(\r_rnd_key_0x[3]_i_58_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[3]_i_53_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[3]_i_54_n_0 ),
        .O(\r_rnd_key_1x[3]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_1x[3]_i_26 
       (.I0(\r_rnd_key_0x[3]_i_55_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[3]_i_56_n_0 ),
        .O(\r_rnd_key_1x[3]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_1x[3]_i_27 
       (.I0(\r_rnd_key_0x[3]_i_65_n_0 ),
        .I1(\r_rnd_key_0x[3]_i_66_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[3]_i_61_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[3]_i_62_n_0 ),
        .O(\r_rnd_key_1x[3]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_1x[3]_i_28 
       (.I0(\r_rnd_key_0x[3]_i_63_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[3]_i_64_n_0 ),
        .O(\r_rnd_key_1x[3]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_1x[3]_i_4 
       (.I0(i_mk[11]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[107]),
        .O(\r_rnd_key_1x[3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_1x[4]_i_1 
       (.I0(w_sk2x_tmp[4]),
        .I1(i_op),
        .I2(w_sk1x_tmp[4]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_1x[4]_i_2_n_0 ),
        .O(\r_rnd_key_1x[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_1x[4]_i_2 
       (.I0(i_mk[12]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[108]),
        .O(\r_rnd_key_1x[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_1x[5]_i_1 
       (.I0(w_sk2x_tmp[5]),
        .I1(i_op),
        .I2(w_sk1x_tmp[5]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_1x[5]_i_2_n_0 ),
        .O(\r_rnd_key_1x[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_1x[5]_i_2 
       (.I0(i_mk[13]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[109]),
        .O(\r_rnd_key_1x[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_1x[6]_i_1 
       (.I0(w_sk2x_tmp[6]),
        .I1(i_op),
        .I2(w_sk1x_tmp[6]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_1x[6]_i_2_n_0 ),
        .O(\r_rnd_key_1x[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_1x[6]_i_2 
       (.I0(i_mk[14]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[110]),
        .O(\r_rnd_key_1x[6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_1x[7]_i_1 
       (.I0(w_sk2x_tmp[7]),
        .I1(i_op),
        .I2(w_sk1x_tmp[7]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_1x[7]_i_4_n_0 ),
        .O(\r_rnd_key_1x[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_1x[7]_i_13 
       (.I0(\r_rnd_key_0x[7]_i_53_n_0 ),
        .I1(\r_rnd_key_0x[7]_i_48_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[7]_i_49_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[7]_i_50_n_0 ),
        .O(\r_rnd_key_1x[7]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_1x[7]_i_14 
       (.I0(\r_rnd_key_0x[7]_i_55_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_52_n_0 ),
        .O(\r_rnd_key_1x[7]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_1x[7]_i_15 
       (.I0(\r_rnd_key_0x[7]_i_61_n_0 ),
        .I1(\r_rnd_key_0x[7]_i_56_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[7]_i_57_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[7]_i_58_n_0 ),
        .O(\r_rnd_key_1x[7]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_1x[7]_i_16 
       (.I0(\r_rnd_key_0x[7]_i_63_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_60_n_0 ),
        .O(\r_rnd_key_1x[7]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_1x[7]_i_17 
       (.I0(\r_rnd_key_0x[7]_i_69_n_0 ),
        .I1(\r_rnd_key_0x[7]_i_64_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[7]_i_65_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[7]_i_66_n_0 ),
        .O(\r_rnd_key_1x[7]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_1x[7]_i_18 
       (.I0(\r_rnd_key_0x[7]_i_71_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_68_n_0 ),
        .O(\r_rnd_key_1x[7]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_1x[7]_i_19 
       (.I0(\r_rnd_key_0x[7]_i_52_n_0 ),
        .I1(\r_rnd_key_0x[7]_i_53_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[7]_i_48_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[7]_i_49_n_0 ),
        .O(\r_rnd_key_1x[7]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_1x[7]_i_20 
       (.I0(\r_rnd_key_0x[7]_i_50_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_51_n_0 ),
        .O(\r_rnd_key_1x[7]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_1x[7]_i_21 
       (.I0(\r_rnd_key_0x[7]_i_60_n_0 ),
        .I1(\r_rnd_key_0x[7]_i_61_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[7]_i_56_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[7]_i_57_n_0 ),
        .O(\r_rnd_key_1x[7]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_1x[7]_i_22 
       (.I0(\r_rnd_key_0x[7]_i_58_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_59_n_0 ),
        .O(\r_rnd_key_1x[7]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_1x[7]_i_23 
       (.I0(\r_rnd_key_0x[7]_i_68_n_0 ),
        .I1(\r_rnd_key_0x[7]_i_69_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I3(\r_rnd_key_0x[7]_i_64_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [2]),
        .I5(\r_rnd_key_0x[7]_i_65_n_0 ),
        .O(\r_rnd_key_1x[7]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_1x[7]_i_24 
       (.I0(\r_rnd_key_0x[7]_i_66_n_0 ),
        .I1(i_op),
        .I2(w_rnd_idx[2]),
        .I3(\r_rnd_key_0x[7]_i_67_n_0 ),
        .O(\r_rnd_key_1x[7]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_1x[7]_i_4 
       (.I0(i_mk[15]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[111]),
        .O(\r_rnd_key_1x[7]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_1x[7]_i_5 
       (.I0(\r_rnd_key_0x[7]_i_28_n_0 ),
        .I1(\r_rnd_key_0x[7]_i_29_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[7]_i_30_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[7]_i_27_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/w_mk2x ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rnd_key_1x[7]_i_9 
       (.I0(\r_rnd_key_0x[7]_i_17_n_0 ),
        .I1(\r_rnd_key_0x[7]_i_14_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[7]_i_15_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[7]_i_16_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/w_mk1x ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_rnd_key_1x_reg[3]_i_2 
       (.CI(\<const0>__0__0 ),
        .CO(r_rnd_key_1x_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({g0_b5_n_0,g0_b4_n_0,g0_b0__0_n_0,g0_b2_n_0}),
        .O(w_sk2x_tmp[3:0]),
        .S({\u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_5_n_0 ,\u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_6_n_0 ,\u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_7_n_0 ,\u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_8_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_rnd_key_1x_reg[3]_i_3 
       (.CI(\<const0>__0__0 ),
        .CO({\r_rnd_key_1x_reg[3]_i_3_n_0 ,\r_rnd_key_1x_reg[3]_i_3_n_1 ,\r_rnd_key_1x_reg[3]_i_3_n_2 ,\r_rnd_key_1x_reg[3]_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({g0_b4_n_0,g0_b0__0_n_0,g0_b2_n_0,g0_b1_n_0}),
        .O(w_sk1x_tmp[3:0]),
        .S({\u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_9_n_0 ,\u_KEY_SCHED/u_SKG/r_rnd_key_1x ,\u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_11_n_0 ,\u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_12_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_rnd_key_1x_reg[7]_i_2 
       (.CI(r_rnd_key_1x_reg[3]),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,g0_b5__0_n_0,g0_b4__0_n_0,g0_b6_n_0}),
        .O(w_sk2x_tmp[7:4]),
        .S({\u_KEY_SCHED/u_SKG/w_mk2x ,\u_KEY_SCHED/u_SKG/r_rnd_key_1x[7]_i_6_n_0 ,\u_KEY_SCHED/u_SKG/r_rnd_key_1x[7]_i_7_n_0 ,\u_KEY_SCHED/u_SKG/r_rnd_key_1x[7]_i_8_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_rnd_key_1x_reg[7]_i_3 
       (.CI(\r_rnd_key_1x_reg[3]_i_3_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,g0_b4__0_n_0,g0_b6_n_0,g0_b5_n_0}),
        .O(w_sk1x_tmp[7:4]),
        .S({\u_KEY_SCHED/u_SKG/w_mk1x ,\u_KEY_SCHED/u_SKG/r_rnd_key_1x[7]_i_10_n_0 ,\u_KEY_SCHED/u_SKG/r_rnd_key_1x[7]_i_11_n_0 ,\u_KEY_SCHED/u_SKG/r_rnd_key_1x[7]_i_12_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_2x[0]_i_1 
       (.I0(w_sk1x_tmp[0]),
        .I1(i_op),
        .I2(w_sk2x_tmp[0]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_2x[0]_i_2_n_0 ),
        .O(r_rnd_key_2x));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_2x[0]_i_2 
       (.I0(i_mk[16]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[112]),
        .O(\r_rnd_key_2x[0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_2x[1]_i_1 
       (.I0(w_sk1x_tmp[1]),
        .I1(i_op),
        .I2(w_sk2x_tmp[1]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_2x[1]_i_2_n_0 ),
        .O(\r_rnd_key_2x[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_2x[1]_i_2 
       (.I0(i_mk[17]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[113]),
        .O(\r_rnd_key_2x[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_2x[2]_i_1 
       (.I0(w_sk1x_tmp[2]),
        .I1(i_op),
        .I2(w_sk2x_tmp[2]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_2x[2]_i_2_n_0 ),
        .O(\r_rnd_key_2x[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_2x[2]_i_2 
       (.I0(i_mk[18]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[114]),
        .O(\r_rnd_key_2x[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_2x[3]_i_1 
       (.I0(w_sk1x_tmp[3]),
        .I1(i_op),
        .I2(w_sk2x_tmp[3]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_2x[3]_i_2_n_0 ),
        .O(\r_rnd_key_2x[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_2x[3]_i_2 
       (.I0(i_mk[19]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[115]),
        .O(\r_rnd_key_2x[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_2x[4]_i_1 
       (.I0(w_sk1x_tmp[4]),
        .I1(i_op),
        .I2(w_sk2x_tmp[4]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_2x[4]_i_2_n_0 ),
        .O(\r_rnd_key_2x[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_2x[4]_i_2 
       (.I0(i_mk[20]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[116]),
        .O(\r_rnd_key_2x[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_2x[5]_i_1 
       (.I0(w_sk1x_tmp[5]),
        .I1(i_op),
        .I2(w_sk2x_tmp[5]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_2x[5]_i_2_n_0 ),
        .O(\r_rnd_key_2x[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_2x[5]_i_2 
       (.I0(i_mk[21]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[117]),
        .O(\r_rnd_key_2x[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_2x[6]_i_1 
       (.I0(w_sk1x_tmp[6]),
        .I1(i_op),
        .I2(w_sk2x_tmp[6]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_2x[6]_i_2_n_0 ),
        .O(\r_rnd_key_2x[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_2x[6]_i_2 
       (.I0(i_mk[22]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[118]),
        .O(\r_rnd_key_2x[6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_2x[7]_i_1 
       (.I0(w_sk1x_tmp[7]),
        .I1(i_op),
        .I2(w_sk2x_tmp[7]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_2x[7]_i_2_n_0 ),
        .O(\r_rnd_key_2x[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_2x[7]_i_2 
       (.I0(i_mk[23]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[119]),
        .O(\r_rnd_key_2x[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_3x[0]_i_1 
       (.I0(w_sk0x_tmp[0]),
        .I1(i_op),
        .I2(w_sk3x_tmp[0]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_3x[0]_i_2_n_0 ),
        .O(r_rnd_key_3x));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_3x[0]_i_2 
       (.I0(i_mk[24]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[120]),
        .O(\r_rnd_key_3x[0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_3x[1]_i_1 
       (.I0(w_sk0x_tmp[1]),
        .I1(i_op),
        .I2(w_sk3x_tmp[1]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_3x[1]_i_2_n_0 ),
        .O(\r_rnd_key_3x[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_3x[1]_i_2 
       (.I0(i_mk[25]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[121]),
        .O(\r_rnd_key_3x[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_3x[2]_i_1 
       (.I0(w_sk0x_tmp[2]),
        .I1(i_op),
        .I2(w_sk3x_tmp[2]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_3x[2]_i_2_n_0 ),
        .O(\r_rnd_key_3x[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_3x[2]_i_2 
       (.I0(i_mk[26]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[122]),
        .O(\r_rnd_key_3x[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_3x[3]_i_1 
       (.I0(w_sk0x_tmp[3]),
        .I1(i_op),
        .I2(w_sk3x_tmp[3]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_3x[3]_i_2_n_0 ),
        .O(\r_rnd_key_3x[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_3x[3]_i_2 
       (.I0(i_mk[27]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[123]),
        .O(\r_rnd_key_3x[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_3x[4]_i_1 
       (.I0(w_sk0x_tmp[4]),
        .I1(i_op),
        .I2(w_sk3x_tmp[4]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_3x[4]_i_2_n_0 ),
        .O(\r_rnd_key_3x[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_3x[4]_i_2 
       (.I0(i_mk[28]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[124]),
        .O(\r_rnd_key_3x[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_3x[5]_i_1 
       (.I0(w_sk0x_tmp[5]),
        .I1(i_op),
        .I2(w_sk3x_tmp[5]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_3x[5]_i_2_n_0 ),
        .O(\r_rnd_key_3x[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_3x[5]_i_2 
       (.I0(i_mk[29]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[125]),
        .O(\r_rnd_key_3x[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_3x[6]_i_1 
       (.I0(w_sk0x_tmp[6]),
        .I1(i_op),
        .I2(w_sk3x_tmp[6]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_3x[6]_i_2_n_0 ),
        .O(\r_rnd_key_3x[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_3x[6]_i_2 
       (.I0(i_mk[30]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[126]),
        .O(\r_rnd_key_3x[6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_rnd_key_3x[7]_i_1 
       (.I0(w_sk0x_tmp[7]),
        .I1(i_op),
        .I2(w_sk3x_tmp[7]),
        .I3(\r_rnd_key_0x[7]_i_4_n_0 ),
        .I4(\r_rnd_key_3x[7]_i_2_n_0 ),
        .O(\r_rnd_key_3x[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEB28)) 
    \r_rnd_key_3x[7]_i_2 
       (.I0(i_mk[31]),
        .I1(w_wf_post_pre),
        .I2(i_op),
        .I3(i_mk[127]),
        .O(\r_rnd_key_3x[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair25" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[0]_i_1 
       (.I0(r_xf),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(\r_xf_reg[3]_i_3_n_7 ),
        .O(p_1_in[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBB88888BB88BB8)) 
    \r_xf[0]_i_2 
       (.I0(o_text_out[0]),
        .I1(w_wf_post_pre),
        .I2(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]15_out [0]),
        .I3(o_text_out[56]),
        .I4(\w_rf_mv[0]0 [0]),
        .I5(i_op),
        .O(r_xf));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[10]_i_1 
       (.I0(\r_xf[10]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[10]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[10]),
        .O(p_1_in[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \r_xf[10]_i_2 
       (.I0(\w_rf_mv[0]00_in [2]),
        .I1(\w_rf_mv[0]0 [2]),
        .I2(w_wf_post_pre),
        .I3(o_text_out[18]),
        .I4(i_op),
        .I5(o_text_out[2]),
        .O(\r_xf[10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[11]_i_1 
       (.I0(\r_xf[11]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[11]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[11]),
        .O(p_1_in[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \r_xf[11]_i_2 
       (.I0(\w_rf_mv[0]00_in [3]),
        .I1(\w_rf_mv[0]0 [3]),
        .I2(w_wf_post_pre),
        .I3(o_text_out[19]),
        .I4(i_op),
        .I5(o_text_out[3]),
        .O(\r_xf[11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[12]_i_1 
       (.I0(\r_xf[12]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[12]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[12]),
        .O(p_1_in[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \r_xf[12]_i_2 
       (.I0(\w_rf_mv[0]00_in [4]),
        .I1(\w_rf_mv[0]0 [4]),
        .I2(w_wf_post_pre),
        .I3(o_text_out[20]),
        .I4(i_op),
        .I5(o_text_out[4]),
        .O(\r_xf[12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[13]_i_1 
       (.I0(\r_xf[13]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[13]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[13]),
        .O(p_1_in[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \r_xf[13]_i_2 
       (.I0(\w_rf_mv[0]00_in [5]),
        .I1(\w_rf_mv[0]0 [5]),
        .I2(w_wf_post_pre),
        .I3(o_text_out[21]),
        .I4(i_op),
        .I5(o_text_out[5]),
        .O(\r_xf[13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[14]_i_1 
       (.I0(\r_xf[14]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[14]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[14]),
        .O(p_1_in[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \r_xf[14]_i_2 
       (.I0(\w_rf_mv[0]00_in [6]),
        .I1(\w_rf_mv[0]0 [6]),
        .I2(w_wf_post_pre),
        .I3(o_text_out[22]),
        .I4(i_op),
        .I5(o_text_out[6]),
        .O(\r_xf[14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[15]_i_1 
       (.I0(\r_xf[15]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[15]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[15]),
        .O(p_1_in[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \r_xf[15]_i_2 
       (.I0(\w_rf_mv[0]00_in [7]),
        .I1(\w_rf_mv[0]0 [7]),
        .I2(w_wf_post_pre),
        .I3(o_text_out[23]),
        .I4(i_op),
        .I5(o_text_out[7]),
        .O(\r_xf[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8B8B8BB8B8B88BB8)) 
    \r_xf[16]_i_1 
       (.I0(\r_xf[16]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(w_rnd_key[8]),
        .I3(i_text_in[16]),
        .I4(\r_xf[55]_i_3_n_0 ),
        .I5(o_text_out[16]),
        .O(p_1_in[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8BBBB8BB88888)) 
    \r_xf[16]_i_2 
       (.I0(o_text_out[16]),
        .I1(w_wf_post_pre),
        .I2(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__43 [0]),
        .I3(o_text_out[24]),
        .I4(i_op),
        .I5(\w_rf_mv[0]00_in [0]),
        .O(\r_xf[16]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8B8B8BB8B8B88BB8)) 
    \r_xf[17]_i_1 
       (.I0(\r_xf[17]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(w_rnd_key[9]),
        .I3(i_text_in[17]),
        .I4(\r_xf[55]_i_3_n_0 ),
        .I5(o_text_out[17]),
        .O(p_1_in[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8BBBB8BB88888)) 
    \r_xf[17]_i_2 
       (.I0(o_text_out[17]),
        .I1(w_wf_post_pre),
        .I2(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__43 [1]),
        .I3(o_text_out[25]),
        .I4(i_op),
        .I5(\w_rf_mv[0]00_in [1]),
        .O(\r_xf[17]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8B8B8BB8B8B88BB8)) 
    \r_xf[18]_i_1 
       (.I0(\r_xf[18]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(w_rnd_key[10]),
        .I3(i_text_in[18]),
        .I4(\r_xf[55]_i_3_n_0 ),
        .I5(o_text_out[18]),
        .O(p_1_in[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8BBBB8BB88888)) 
    \r_xf[18]_i_2 
       (.I0(o_text_out[18]),
        .I1(w_wf_post_pre),
        .I2(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__43 [2]),
        .I3(o_text_out[26]),
        .I4(i_op),
        .I5(\w_rf_mv[0]00_in [2]),
        .O(\r_xf[18]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8B8B8BB8B8B88BB8)) 
    \r_xf[19]_i_1 
       (.I0(\r_xf[19]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(w_rnd_key[11]),
        .I3(i_text_in[19]),
        .I4(\r_xf[55]_i_3_n_0 ),
        .I5(o_text_out[19]),
        .O(p_1_in[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8BBBB8BB88888)) 
    \r_xf[19]_i_2 
       (.I0(o_text_out[19]),
        .I1(w_wf_post_pre),
        .I2(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__43 [3]),
        .I3(o_text_out[27]),
        .I4(i_op),
        .I5(\w_rf_mv[0]00_in [3]),
        .O(\r_xf[19]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair25" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[1]_i_1 
       (.I0(\r_xf[1]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(\r_xf_reg[3]_i_3_n_6 ),
        .O(p_1_in[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBB88888BB88BB8)) 
    \r_xf[1]_i_2 
       (.I0(o_text_out[1]),
        .I1(w_wf_post_pre),
        .I2(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]15_out [1]),
        .I3(o_text_out[57]),
        .I4(\w_rf_mv[0]0 [1]),
        .I5(i_op),
        .O(\r_xf[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8B8B8BB8B8B88BB8)) 
    \r_xf[20]_i_1 
       (.I0(\r_xf[20]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(w_rnd_key[12]),
        .I3(i_text_in[20]),
        .I4(\r_xf[55]_i_3_n_0 ),
        .I5(o_text_out[20]),
        .O(p_1_in[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8BBBB8BB88888)) 
    \r_xf[20]_i_2 
       (.I0(o_text_out[20]),
        .I1(w_wf_post_pre),
        .I2(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__43 [4]),
        .I3(o_text_out[28]),
        .I4(i_op),
        .I5(\w_rf_mv[0]00_in [4]),
        .O(\r_xf[20]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8B8B8BB8B8B88BB8)) 
    \r_xf[21]_i_1 
       (.I0(\r_xf[21]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(w_rnd_key[13]),
        .I3(i_text_in[21]),
        .I4(\r_xf[55]_i_3_n_0 ),
        .I5(o_text_out[21]),
        .O(p_1_in[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8BBBB8BB88888)) 
    \r_xf[21]_i_2 
       (.I0(o_text_out[21]),
        .I1(w_wf_post_pre),
        .I2(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__43 [5]),
        .I3(o_text_out[29]),
        .I4(i_op),
        .I5(\w_rf_mv[0]00_in [5]),
        .O(\r_xf[21]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8B8B8BB8B8B88BB8)) 
    \r_xf[22]_i_1 
       (.I0(\r_xf[22]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(w_rnd_key[14]),
        .I3(i_text_in[22]),
        .I4(\r_xf[55]_i_3_n_0 ),
        .I5(o_text_out[22]),
        .O(p_1_in[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8BBBB8BB88888)) 
    \r_xf[22]_i_2 
       (.I0(o_text_out[22]),
        .I1(w_wf_post_pre),
        .I2(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__43 [6]),
        .I3(o_text_out[30]),
        .I4(i_op),
        .I5(\w_rf_mv[0]00_in [6]),
        .O(\r_xf[22]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8B8B8BB8B8B88BB8)) 
    \r_xf[23]_i_1 
       (.I0(\r_xf[23]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(w_rnd_key[15]),
        .I3(i_text_in[23]),
        .I4(\r_xf[55]_i_3_n_0 ),
        .I5(o_text_out[23]),
        .O(p_1_in[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8BBBB8BB88888)) 
    \r_xf[23]_i_2 
       (.I0(o_text_out[23]),
        .I1(w_wf_post_pre),
        .I2(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__43 [7]),
        .I3(o_text_out[31]),
        .I4(i_op),
        .I5(\w_rf_mv[0]00_in [7]),
        .O(\r_xf[23]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[24]_i_1 
       (.I0(\r_xf[24]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[24]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[24]),
        .O(p_1_in[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1DE2FFFF1DE20000)) 
    \r_xf[24]_i_2 
       (.I0(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]12_out [0]),
        .I1(i_op),
        .I2(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__43 [0]),
        .I3(o_text_out[24]),
        .I4(w_wf_post_pre),
        .I5(\r_xf[24]_i_3_n_0 ),
        .O(\r_xf[24]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[24]_i_3 
       (.I0(o_text_out[32]),
        .I1(i_op),
        .I2(o_text_out[16]),
        .O(\r_xf[24]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[25]_i_1 
       (.I0(\r_xf[25]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[25]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[25]),
        .O(p_1_in[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1DE2FFFF1DE20000)) 
    \r_xf[25]_i_2 
       (.I0(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]12_out [1]),
        .I1(i_op),
        .I2(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__43 [1]),
        .I3(o_text_out[25]),
        .I4(w_wf_post_pre),
        .I5(\r_xf[25]_i_3_n_0 ),
        .O(\r_xf[25]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[25]_i_3 
       (.I0(o_text_out[33]),
        .I1(i_op),
        .I2(o_text_out[17]),
        .O(\r_xf[25]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[26]_i_1 
       (.I0(\r_xf[26]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[26]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[26]),
        .O(p_1_in[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1DE2FFFF1DE20000)) 
    \r_xf[26]_i_2 
       (.I0(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]12_out [2]),
        .I1(i_op),
        .I2(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__43 [2]),
        .I3(o_text_out[26]),
        .I4(w_wf_post_pre),
        .I5(\r_xf[26]_i_3_n_0 ),
        .O(\r_xf[26]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[26]_i_3 
       (.I0(o_text_out[34]),
        .I1(i_op),
        .I2(o_text_out[18]),
        .O(\r_xf[26]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[27]_i_1 
       (.I0(\r_xf[27]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[27]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[27]),
        .O(p_1_in[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1DE2FFFF1DE20000)) 
    \r_xf[27]_i_2 
       (.I0(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]12_out [3]),
        .I1(i_op),
        .I2(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__43 [3]),
        .I3(o_text_out[27]),
        .I4(w_wf_post_pre),
        .I5(\r_xf[27]_i_3_n_0 ),
        .O(\r_xf[27]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[27]_i_3 
       (.I0(o_text_out[35]),
        .I1(i_op),
        .I2(o_text_out[19]),
        .O(\r_xf[27]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[28]_i_1 
       (.I0(\r_xf[28]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[28]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[28]),
        .O(p_1_in[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1DE2FFFF1DE20000)) 
    \r_xf[28]_i_2 
       (.I0(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]12_out [4]),
        .I1(i_op),
        .I2(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__43 [4]),
        .I3(o_text_out[28]),
        .I4(w_wf_post_pre),
        .I5(\r_xf[28]_i_3_n_0 ),
        .O(\r_xf[28]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[28]_i_3 
       (.I0(o_text_out[36]),
        .I1(i_op),
        .I2(o_text_out[20]),
        .O(\r_xf[28]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[29]_i_1 
       (.I0(\r_xf[29]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[29]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[29]),
        .O(p_1_in[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1DE2FFFF1DE20000)) 
    \r_xf[29]_i_2 
       (.I0(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]12_out [5]),
        .I1(i_op),
        .I2(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__43 [5]),
        .I3(o_text_out[29]),
        .I4(w_wf_post_pre),
        .I5(\r_xf[29]_i_3_n_0 ),
        .O(\r_xf[29]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[29]_i_3 
       (.I0(o_text_out[37]),
        .I1(i_op),
        .I2(o_text_out[21]),
        .O(\r_xf[29]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair26" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[2]_i_1 
       (.I0(\r_xf[2]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(\r_xf_reg[3]_i_3_n_5 ),
        .O(p_1_in[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBB88888BB88BB8)) 
    \r_xf[2]_i_2 
       (.I0(o_text_out[2]),
        .I1(w_wf_post_pre),
        .I2(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]15_out [2]),
        .I3(o_text_out[58]),
        .I4(\w_rf_mv[0]0 [2]),
        .I5(i_op),
        .O(\r_xf[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[30]_i_1 
       (.I0(\r_xf[30]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[30]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[30]),
        .O(p_1_in[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1DE2FFFF1DE20000)) 
    \r_xf[30]_i_2 
       (.I0(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]12_out [6]),
        .I1(i_op),
        .I2(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__43 [6]),
        .I3(o_text_out[30]),
        .I4(w_wf_post_pre),
        .I5(\r_xf[30]_i_3_n_0 ),
        .O(\r_xf[30]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[30]_i_3 
       (.I0(o_text_out[38]),
        .I1(i_op),
        .I2(o_text_out[22]),
        .O(\r_xf[30]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[31]_i_1 
       (.I0(\r_xf[31]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[31]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[31]),
        .O(p_1_in[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1DE2FFFF1DE20000)) 
    \r_xf[31]_i_2 
       (.I0(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]12_out [7]),
        .I1(i_op),
        .I2(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__43 [7]),
        .I3(o_text_out[31]),
        .I4(w_wf_post_pre),
        .I5(\r_xf[31]_i_3_n_0 ),
        .O(\r_xf[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[31]_i_3 
       (.I0(o_text_out[39]),
        .I1(i_op),
        .I2(o_text_out[23]),
        .O(\r_xf[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair29" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[32]_i_1 
       (.I0(\r_xf[32]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(\r_xf_reg[35]_i_3_n_7 ),
        .O(p_1_in[32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888B8BBB8BBB888)) 
    \r_xf[32]_i_2 
       (.I0(o_text_out[32]),
        .I1(w_wf_post_pre),
        .I2(\w_rf_mv[2]0 [0]),
        .I3(i_op),
        .I4(o_text_out[24]),
        .I5(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]12_out [0]),
        .O(\r_xf[32]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair32" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[33]_i_1 
       (.I0(\r_xf[33]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(\r_xf_reg[35]_i_3_n_6 ),
        .O(p_1_in[33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888B8BBB8BBB888)) 
    \r_xf[33]_i_2 
       (.I0(o_text_out[33]),
        .I1(w_wf_post_pre),
        .I2(\w_rf_mv[2]0 [1]),
        .I3(i_op),
        .I4(o_text_out[25]),
        .I5(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]12_out [1]),
        .O(\r_xf[33]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair32" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[34]_i_1 
       (.I0(\r_xf[34]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(\r_xf_reg[35]_i_3_n_5 ),
        .O(p_1_in[34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888B8BBB8BBB888)) 
    \r_xf[34]_i_2 
       (.I0(o_text_out[34]),
        .I1(w_wf_post_pre),
        .I2(\w_rf_mv[2]0 [2]),
        .I3(i_op),
        .I4(o_text_out[26]),
        .I5(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]12_out [2]),
        .O(\r_xf[34]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair35" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[35]_i_1 
       (.I0(\r_xf[35]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(\r_xf_reg[35]_i_3_n_4 ),
        .O(p_1_in[35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9699999996666666)) 
    \r_xf[35]_i_10 
       (.I0(w_rnd_key[17]),
        .I1(i_op),
        .I2(i_text_in[33]),
        .I3(i_text_val),
        .I4(o_rdy_INST_0_i_1_n_0),
        .I5(o_text_out[33]),
        .O(\r_xf[35]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888B8BBB8BBB888)) 
    \r_xf[35]_i_2 
       (.I0(o_text_out[35]),
        .I1(w_wf_post_pre),
        .I2(\w_rf_mv[2]0 [3]),
        .I3(i_op),
        .I4(o_text_out[27]),
        .I5(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]12_out [3]),
        .O(\r_xf[35]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEA2A)) 
    \r_xf[35]_i_4 
       (.I0(o_text_out[32]),
        .I1(o_rdy_INST_0_i_1_n_0),
        .I2(i_text_val),
        .I3(i_text_in[32]),
        .O(\u_CRYPTO_PATH/w_wf_in_mux [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_xf[35]_i_5 
       (.I0(i_op),
        .I1(w_rnd_key[19]),
        .O(\r_xf[35]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_xf[35]_i_6 
       (.I0(i_op),
        .I1(w_rnd_key[18]),
        .O(\r_xf[35]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_xf[35]_i_7 
       (.I0(i_op),
        .I1(w_rnd_key[17]),
        .O(\r_xf[35]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9699999996666666)) 
    \r_xf[35]_i_8 
       (.I0(w_rnd_key[19]),
        .I1(i_op),
        .I2(i_text_in[35]),
        .I3(i_text_val),
        .I4(o_rdy_INST_0_i_1_n_0),
        .I5(o_text_out[35]),
        .O(\r_xf[35]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9699999996666666)) 
    \r_xf[35]_i_9 
       (.I0(w_rnd_key[18]),
        .I1(i_op),
        .I2(i_text_in[34]),
        .I3(i_text_val),
        .I4(o_rdy_INST_0_i_1_n_0),
        .I5(o_text_out[34]),
        .O(\r_xf[35]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair35" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[36]_i_1 
       (.I0(\r_xf[36]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(\r_xf_reg[39]_i_3_n_7 ),
        .O(p_1_in[36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888B8BBB8BBB888)) 
    \r_xf[36]_i_2 
       (.I0(o_text_out[36]),
        .I1(w_wf_post_pre),
        .I2(\w_rf_mv[2]0 [4]),
        .I3(i_op),
        .I4(o_text_out[28]),
        .I5(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]12_out [4]),
        .O(\r_xf[36]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair38" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[37]_i_1 
       (.I0(\r_xf[37]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(\r_xf_reg[39]_i_3_n_6 ),
        .O(p_1_in[37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888B8BBB8BBB888)) 
    \r_xf[37]_i_2 
       (.I0(o_text_out[37]),
        .I1(w_wf_post_pre),
        .I2(\w_rf_mv[2]0 [5]),
        .I3(i_op),
        .I4(o_text_out[29]),
        .I5(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]12_out [5]),
        .O(\r_xf[37]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair38" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[38]_i_1 
       (.I0(\r_xf[38]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(\r_xf_reg[39]_i_3_n_5 ),
        .O(p_1_in[38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888B8BBB8BBB888)) 
    \r_xf[38]_i_2 
       (.I0(o_text_out[38]),
        .I1(w_wf_post_pre),
        .I2(\w_rf_mv[2]0 [6]),
        .I3(i_op),
        .I4(o_text_out[30]),
        .I5(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]12_out [6]),
        .O(\r_xf[38]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair27" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[39]_i_1 
       (.I0(\r_xf[39]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(\r_xf_reg[39]_i_3_n_4 ),
        .O(p_1_in[39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9699999996666666)) 
    \r_xf[39]_i_10 
       (.I0(w_rnd_key[20]),
        .I1(i_op),
        .I2(i_text_in[36]),
        .I3(i_text_val),
        .I4(o_rdy_INST_0_i_1_n_0),
        .I5(o_text_out[36]),
        .O(\r_xf[39]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888B8BBB8BBB888)) 
    \r_xf[39]_i_2 
       (.I0(o_text_out[39]),
        .I1(w_wf_post_pre),
        .I2(\w_rf_mv[2]0 [7]),
        .I3(i_op),
        .I4(o_text_out[31]),
        .I5(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]12_out [7]),
        .O(\r_xf[39]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_xf[39]_i_4 
       (.I0(i_op),
        .I1(w_rnd_key[22]),
        .O(\r_xf[39]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_xf[39]_i_5 
       (.I0(i_op),
        .I1(w_rnd_key[21]),
        .O(\r_xf[39]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_xf[39]_i_6 
       (.I0(i_op),
        .I1(w_rnd_key[20]),
        .O(\r_xf[39]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBF80407F407FBF80)) 
    \r_xf[39]_i_7 
       (.I0(i_text_in[39]),
        .I1(i_text_val),
        .I2(o_rdy_INST_0_i_1_n_0),
        .I3(o_text_out[39]),
        .I4(w_rnd_key[23]),
        .I5(i_op),
        .O(\r_xf[39]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9699999996666666)) 
    \r_xf[39]_i_8 
       (.I0(w_rnd_key[22]),
        .I1(i_op),
        .I2(i_text_in[38]),
        .I3(i_text_val),
        .I4(o_rdy_INST_0_i_1_n_0),
        .I5(o_text_out[38]),
        .O(\r_xf[39]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9699999996666666)) 
    \r_xf[39]_i_9 
       (.I0(w_rnd_key[21]),
        .I1(i_op),
        .I2(i_text_in[37]),
        .I3(i_text_val),
        .I4(o_rdy_INST_0_i_1_n_0),
        .I5(o_text_out[37]),
        .O(\r_xf[39]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair26" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[3]_i_1 
       (.I0(\r_xf[3]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(\r_xf_reg[3]_i_3_n_4 ),
        .O(p_1_in[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9699999996666666)) 
    \r_xf[3]_i_10 
       (.I0(w_rnd_key[1]),
        .I1(i_op),
        .I2(i_text_in[1]),
        .I3(i_text_val),
        .I4(o_rdy_INST_0_i_1_n_0),
        .I5(o_text_out[1]),
        .O(\r_xf[3]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBB88888BB88BB8)) 
    \r_xf[3]_i_2 
       (.I0(o_text_out[3]),
        .I1(w_wf_post_pre),
        .I2(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]15_out [3]),
        .I3(o_text_out[59]),
        .I4(\w_rf_mv[0]0 [3]),
        .I5(i_op),
        .O(\r_xf[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEA2A)) 
    \r_xf[3]_i_4 
       (.I0(o_text_out[0]),
        .I1(o_rdy_INST_0_i_1_n_0),
        .I2(i_text_val),
        .I3(i_text_in[0]),
        .O(\u_CRYPTO_PATH/w_wf_in_mux [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_xf[3]_i_5 
       (.I0(i_op),
        .I1(w_rnd_key[3]),
        .O(\r_xf[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_xf[3]_i_6 
       (.I0(i_op),
        .I1(w_rnd_key[2]),
        .O(\r_xf[3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_xf[3]_i_7 
       (.I0(i_op),
        .I1(w_rnd_key[1]),
        .O(\r_xf[3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9699999996666666)) 
    \r_xf[3]_i_8 
       (.I0(w_rnd_key[3]),
        .I1(i_op),
        .I2(i_text_in[3]),
        .I3(i_text_val),
        .I4(o_rdy_INST_0_i_1_n_0),
        .I5(o_text_out[3]),
        .O(\r_xf[3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9699999996666666)) 
    \r_xf[3]_i_9 
       (.I0(w_rnd_key[2]),
        .I1(i_op),
        .I2(i_text_in[2]),
        .I3(i_text_val),
        .I4(o_rdy_INST_0_i_1_n_0),
        .I5(o_text_out[2]),
        .O(\r_xf[3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[40]_i_1 
       (.I0(\r_xf[40]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[40]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[40]),
        .O(p_1_in[40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \r_xf[40]_i_2 
       (.I0(\w_rf_mv[2]01_in [0]),
        .I1(\w_rf_mv[2]0 [0]),
        .I2(w_wf_post_pre),
        .I3(o_text_out[48]),
        .I4(i_op),
        .I5(o_text_out[32]),
        .O(\r_xf[40]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[41]_i_1 
       (.I0(\r_xf[41]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[41]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[41]),
        .O(p_1_in[41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \r_xf[41]_i_2 
       (.I0(\w_rf_mv[2]01_in [1]),
        .I1(\w_rf_mv[2]0 [1]),
        .I2(w_wf_post_pre),
        .I3(o_text_out[49]),
        .I4(i_op),
        .I5(o_text_out[33]),
        .O(\r_xf[41]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[42]_i_1 
       (.I0(\r_xf[42]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[42]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[42]),
        .O(p_1_in[42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \r_xf[42]_i_2 
       (.I0(\w_rf_mv[2]01_in [2]),
        .I1(\w_rf_mv[2]0 [2]),
        .I2(w_wf_post_pre),
        .I3(o_text_out[50]),
        .I4(i_op),
        .I5(o_text_out[34]),
        .O(\r_xf[42]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[43]_i_1 
       (.I0(\r_xf[43]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[43]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[43]),
        .O(p_1_in[43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \r_xf[43]_i_2 
       (.I0(\w_rf_mv[2]01_in [3]),
        .I1(\w_rf_mv[2]0 [3]),
        .I2(w_wf_post_pre),
        .I3(o_text_out[51]),
        .I4(i_op),
        .I5(o_text_out[35]),
        .O(\r_xf[43]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[44]_i_1 
       (.I0(\r_xf[44]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[44]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[44]),
        .O(p_1_in[44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \r_xf[44]_i_2 
       (.I0(\w_rf_mv[2]01_in [4]),
        .I1(\w_rf_mv[2]0 [4]),
        .I2(w_wf_post_pre),
        .I3(o_text_out[52]),
        .I4(i_op),
        .I5(o_text_out[36]),
        .O(\r_xf[44]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[45]_i_1 
       (.I0(\r_xf[45]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[45]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[45]),
        .O(p_1_in[45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \r_xf[45]_i_2 
       (.I0(\w_rf_mv[2]01_in [5]),
        .I1(\w_rf_mv[2]0 [5]),
        .I2(w_wf_post_pre),
        .I3(o_text_out[53]),
        .I4(i_op),
        .I5(o_text_out[37]),
        .O(\r_xf[45]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[46]_i_1 
       (.I0(\r_xf[46]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[46]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[46]),
        .O(p_1_in[46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \r_xf[46]_i_2 
       (.I0(\w_rf_mv[2]01_in [6]),
        .I1(\w_rf_mv[2]0 [6]),
        .I2(w_wf_post_pre),
        .I3(o_text_out[54]),
        .I4(i_op),
        .I5(o_text_out[38]),
        .O(\r_xf[46]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[47]_i_1 
       (.I0(\r_xf[47]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[47]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[47]),
        .O(p_1_in[47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \r_xf[47]_i_2 
       (.I0(\w_rf_mv[2]01_in [7]),
        .I1(\w_rf_mv[2]0 [7]),
        .I2(w_wf_post_pre),
        .I3(o_text_out[55]),
        .I4(i_op),
        .I5(o_text_out[39]),
        .O(\r_xf[47]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8B8B8BB8B8B88BB8)) 
    \r_xf[48]_i_1 
       (.I0(\r_xf[48]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(w_rnd_key[24]),
        .I3(i_text_in[48]),
        .I4(\r_xf[55]_i_3_n_0 ),
        .I5(o_text_out[48]),
        .O(p_1_in[48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8BBBB8BB88888)) 
    \r_xf[48]_i_2 
       (.I0(o_text_out[48]),
        .I1(w_wf_post_pre),
        .I2(o_text_out[56]),
        .I3(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__43 [0]),
        .I4(i_op),
        .I5(\w_rf_mv[2]01_in [0]),
        .O(\r_xf[48]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8B8B8BB8B8B88BB8)) 
    \r_xf[49]_i_1 
       (.I0(\r_xf[49]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(w_rnd_key[25]),
        .I3(i_text_in[49]),
        .I4(\r_xf[55]_i_3_n_0 ),
        .I5(o_text_out[49]),
        .O(p_1_in[49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8BBBB8BB88888)) 
    \r_xf[49]_i_2 
       (.I0(o_text_out[49]),
        .I1(w_wf_post_pre),
        .I2(o_text_out[57]),
        .I3(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__43 [1]),
        .I4(i_op),
        .I5(\w_rf_mv[2]01_in [1]),
        .O(\r_xf[49]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair27" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[4]_i_1 
       (.I0(\r_xf[4]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(\r_xf_reg[7]_i_3_n_7 ),
        .O(p_1_in[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBB88888BB88BB8)) 
    \r_xf[4]_i_2 
       (.I0(o_text_out[4]),
        .I1(w_wf_post_pre),
        .I2(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]15_out [4]),
        .I3(o_text_out[60]),
        .I4(\w_rf_mv[0]0 [4]),
        .I5(i_op),
        .O(\r_xf[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8B8B8BB8B8B88BB8)) 
    \r_xf[50]_i_1 
       (.I0(\r_xf[50]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(w_rnd_key[26]),
        .I3(i_text_in[50]),
        .I4(\r_xf[55]_i_3_n_0 ),
        .I5(o_text_out[50]),
        .O(p_1_in[50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8BBBB8BB88888)) 
    \r_xf[50]_i_2 
       (.I0(o_text_out[50]),
        .I1(w_wf_post_pre),
        .I2(o_text_out[58]),
        .I3(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__43 [2]),
        .I4(i_op),
        .I5(\w_rf_mv[2]01_in [2]),
        .O(\r_xf[50]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8B8B8BB8B8B88BB8)) 
    \r_xf[51]_i_1 
       (.I0(\r_xf[51]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(w_rnd_key[27]),
        .I3(i_text_in[51]),
        .I4(\r_xf[55]_i_3_n_0 ),
        .I5(o_text_out[51]),
        .O(p_1_in[51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8BBBB8BB88888)) 
    \r_xf[51]_i_2 
       (.I0(o_text_out[51]),
        .I1(w_wf_post_pre),
        .I2(o_text_out[59]),
        .I3(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__43 [3]),
        .I4(i_op),
        .I5(\w_rf_mv[2]01_in [3]),
        .O(\r_xf[51]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8B8B8BB8B8B88BB8)) 
    \r_xf[52]_i_1 
       (.I0(\r_xf[52]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(w_rnd_key[28]),
        .I3(i_text_in[52]),
        .I4(\r_xf[55]_i_3_n_0 ),
        .I5(o_text_out[52]),
        .O(p_1_in[52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8BBBB8BB88888)) 
    \r_xf[52]_i_2 
       (.I0(o_text_out[52]),
        .I1(w_wf_post_pre),
        .I2(o_text_out[60]),
        .I3(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__43 [4]),
        .I4(i_op),
        .I5(\w_rf_mv[2]01_in [4]),
        .O(\r_xf[52]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8B8B8BB8B8B88BB8)) 
    \r_xf[53]_i_1 
       (.I0(\r_xf[53]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(w_rnd_key[29]),
        .I3(i_text_in[53]),
        .I4(\r_xf[55]_i_3_n_0 ),
        .I5(o_text_out[53]),
        .O(p_1_in[53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8BBBB8BB88888)) 
    \r_xf[53]_i_2 
       (.I0(o_text_out[53]),
        .I1(w_wf_post_pre),
        .I2(o_text_out[61]),
        .I3(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__43 [5]),
        .I4(i_op),
        .I5(\w_rf_mv[2]01_in [5]),
        .O(\r_xf[53]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8B8B8BB8B8B88BB8)) 
    \r_xf[54]_i_1 
       (.I0(\r_xf[54]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(w_rnd_key[30]),
        .I3(i_text_in[54]),
        .I4(\r_xf[55]_i_3_n_0 ),
        .I5(o_text_out[54]),
        .O(p_1_in[54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8BBBB8BB88888)) 
    \r_xf[54]_i_2 
       (.I0(o_text_out[54]),
        .I1(w_wf_post_pre),
        .I2(o_text_out[62]),
        .I3(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__43 [6]),
        .I4(i_op),
        .I5(\w_rf_mv[2]01_in [6]),
        .O(\r_xf[54]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8B8B8BB8B8B88BB8)) 
    \r_xf[55]_i_1 
       (.I0(\r_xf[55]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(w_rnd_key[31]),
        .I3(i_text_in[55]),
        .I4(\r_xf[55]_i_3_n_0 ),
        .I5(o_text_out[55]),
        .O(p_1_in[55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8BBBB8BB88888)) 
    \r_xf[55]_i_2 
       (.I0(o_text_out[55]),
        .I1(w_wf_post_pre),
        .I2(o_text_out[63]),
        .I3(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__43 [7]),
        .I4(i_op),
        .I5(\w_rf_mv[2]01_in [7]),
        .O(\r_xf[55]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \r_xf[55]_i_3 
       (.I0(o_rdy_INST_0_i_1_n_0),
        .I1(i_text_val),
        .O(\r_xf[55]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[56]_i_1 
       (.I0(\r_xf[56]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[56]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[56]),
        .O(p_1_in[56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1ED2FFFF1ED20000)) 
    \r_xf[56]_i_2 
       (.I0(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]15_out [0]),
        .I1(i_op),
        .I2(o_text_out[56]),
        .I3(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__43 [0]),
        .I4(w_wf_post_pre),
        .I5(\r_xf[56]_i_3_n_0 ),
        .O(\r_xf[56]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[56]_i_3 
       (.I0(o_text_out[0]),
        .I1(i_op),
        .I2(o_text_out[48]),
        .O(\r_xf[56]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[57]_i_1 
       (.I0(\r_xf[57]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[57]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[57]),
        .O(p_1_in[57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1ED2FFFF1ED20000)) 
    \r_xf[57]_i_2 
       (.I0(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]15_out [1]),
        .I1(i_op),
        .I2(o_text_out[57]),
        .I3(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__43 [1]),
        .I4(w_wf_post_pre),
        .I5(\r_xf[57]_i_3_n_0 ),
        .O(\r_xf[57]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[57]_i_3 
       (.I0(o_text_out[1]),
        .I1(i_op),
        .I2(o_text_out[49]),
        .O(\r_xf[57]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[58]_i_1 
       (.I0(\r_xf[58]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[58]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[58]),
        .O(p_1_in[58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1ED2FFFF1ED20000)) 
    \r_xf[58]_i_2 
       (.I0(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]15_out [2]),
        .I1(i_op),
        .I2(o_text_out[58]),
        .I3(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__43 [2]),
        .I4(w_wf_post_pre),
        .I5(\r_xf[58]_i_3_n_0 ),
        .O(\r_xf[58]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[58]_i_3 
       (.I0(o_text_out[2]),
        .I1(i_op),
        .I2(o_text_out[50]),
        .O(\r_xf[58]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[59]_i_1 
       (.I0(\r_xf[59]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[59]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[59]),
        .O(p_1_in[59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1ED2FFFF1ED20000)) 
    \r_xf[59]_i_2 
       (.I0(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]15_out [3]),
        .I1(i_op),
        .I2(o_text_out[59]),
        .I3(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__43 [3]),
        .I4(w_wf_post_pre),
        .I5(\r_xf[59]_i_3_n_0 ),
        .O(\r_xf[59]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[59]_i_3 
       (.I0(o_text_out[3]),
        .I1(i_op),
        .I2(o_text_out[51]),
        .O(\r_xf[59]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair28" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[5]_i_1 
       (.I0(\r_xf[5]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(\r_xf_reg[7]_i_3_n_6 ),
        .O(p_1_in[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBB88888BB88BB8)) 
    \r_xf[5]_i_2 
       (.I0(o_text_out[5]),
        .I1(w_wf_post_pre),
        .I2(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]15_out [5]),
        .I3(o_text_out[61]),
        .I4(\w_rf_mv[0]0 [5]),
        .I5(i_op),
        .O(\r_xf[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[60]_i_1 
       (.I0(\r_xf[60]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[60]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[60]),
        .O(p_1_in[60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1ED2FFFF1ED20000)) 
    \r_xf[60]_i_2 
       (.I0(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]15_out [4]),
        .I1(i_op),
        .I2(o_text_out[60]),
        .I3(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__43 [4]),
        .I4(w_wf_post_pre),
        .I5(\r_xf[60]_i_3_n_0 ),
        .O(\r_xf[60]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[60]_i_3 
       (.I0(o_text_out[4]),
        .I1(i_op),
        .I2(o_text_out[52]),
        .O(\r_xf[60]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[61]_i_1 
       (.I0(\r_xf[61]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[61]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[61]),
        .O(p_1_in[61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1ED2FFFF1ED20000)) 
    \r_xf[61]_i_2 
       (.I0(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]15_out [5]),
        .I1(i_op),
        .I2(o_text_out[61]),
        .I3(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__43 [5]),
        .I4(w_wf_post_pre),
        .I5(\r_xf[61]_i_3_n_0 ),
        .O(\r_xf[61]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[61]_i_3 
       (.I0(o_text_out[5]),
        .I1(i_op),
        .I2(o_text_out[53]),
        .O(\r_xf[61]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[62]_i_1 
       (.I0(\r_xf[62]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[62]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[62]),
        .O(p_1_in[62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1ED2FFFF1ED20000)) 
    \r_xf[62]_i_2 
       (.I0(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]15_out [6]),
        .I1(i_op),
        .I2(o_text_out[62]),
        .I3(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__43 [6]),
        .I4(w_wf_post_pre),
        .I5(\r_xf[62]_i_3_n_0 ),
        .O(\r_xf[62]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[62]_i_3 
       (.I0(o_text_out[6]),
        .I1(i_op),
        .I2(o_text_out[54]),
        .O(\r_xf[62]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF2F2F2)) 
    \r_xf[63]_i_1 
       (.I0(\r_xf[63]_i_4_n_0 ),
        .I1(\u_CONTROL/r_pstate_reg ),
        .I2(w_wf_post_pre),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(\u_CONTROL/o_xf_sel2 ),
        .O(\r_xf[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[63]_i_10 
       (.I0(o_text_out[7]),
        .I1(i_op),
        .I2(o_text_out[55]),
        .O(\r_xf[63]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[63]_i_2 
       (.I0(\r_xf[63]_i_8_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[63]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[63]),
        .O(p_1_in[63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \r_xf[63]_i_3 
       (.I0(rstn),
        .O(\r_xf[63]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFD)) 
    \r_xf[63]_i_4 
       (.I0(\u_CONTROL/r_pstate [1]),
        .I1(\u_CONTROL/r_pstate [4]),
        .I2(\u_CONTROL/r_pstate [2]),
        .I3(\u_CONTROL/r_pstate [3]),
        .I4(\u_CONTROL/r_pstate [0]),
        .I5(\u_CONTROL/r_pstate [5]),
        .O(\r_xf[63]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0005000000090009)) 
    \r_xf[63]_i_5 
       (.I0(\u_CONTROL/r_pstate [2]),
        .I1(\u_CONTROL/r_pstate [5]),
        .I2(\u_CONTROL/r_pstate [4]),
        .I3(\u_CONTROL/r_pstate [3]),
        .I4(\u_CONTROL/r_pstate [0]),
        .I5(\u_CONTROL/r_pstate [1]),
        .O(\u_CONTROL/r_pstate_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \r_xf[63]_i_6 
       (.I0(\u_CONTROL/r_pstate [2]),
        .I1(\u_CONTROL/r_pstate [1]),
        .I2(\u_CONTROL/r_pstate [4]),
        .I3(\u_CONTROL/r_pstate [3]),
        .I4(\u_CONTROL/r_pstate [5]),
        .I5(\u_CONTROL/r_pstate [0]),
        .O(w_wf_post_pre));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \r_xf[63]_i_7 
       (.I0(\u_CONTROL/r_pstate [1]),
        .I1(\u_CONTROL/r_pstate [4]),
        .I2(\u_CONTROL/r_pstate [0]),
        .I3(\u_CONTROL/r_pstate [3]),
        .I4(\u_CONTROL/r_pstate [5]),
        .I5(\u_CONTROL/r_pstate [2]),
        .O(\u_CONTROL/o_xf_sel2 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1ED2FFFF1ED20000)) 
    \r_xf[63]_i_8 
       (.I0(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]15_out [7]),
        .I1(i_op),
        .I2(o_text_out[63]),
        .I3(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__43 [7]),
        .I4(w_wf_post_pre),
        .I5(\r_xf[63]_i_10_n_0 ),
        .O(\r_xf[63]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7077707077777777)) 
    \r_xf[63]_i_9 
       (.I0(i_text_val),
        .I1(o_rdy_INST_0_i_1_n_0),
        .I2(w_wf_post_pre),
        .I3(\u_CONTROL/r_pstate_reg ),
        .I4(\r_xf[63]_i_4_n_0 ),
        .I5(\u_CONTROL/o_xf_sel2 ),
        .O(\r_xf[63]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair28" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[6]_i_1 
       (.I0(\r_xf[6]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(\r_xf_reg[7]_i_3_n_5 ),
        .O(p_1_in[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBB88888BB88BB8)) 
    \r_xf[6]_i_2 
       (.I0(o_text_out[6]),
        .I1(w_wf_post_pre),
        .I2(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]15_out [6]),
        .I3(o_text_out[62]),
        .I4(\w_rf_mv[0]0 [6]),
        .I5(i_op),
        .O(\r_xf[6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair29" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_xf[7]_i_1 
       (.I0(\r_xf[7]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(\r_xf_reg[7]_i_3_n_4 ),
        .O(p_1_in[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9699999996666666)) 
    \r_xf[7]_i_10 
       (.I0(w_rnd_key[4]),
        .I1(i_op),
        .I2(i_text_in[4]),
        .I3(i_text_val),
        .I4(o_rdy_INST_0_i_1_n_0),
        .I5(o_text_out[4]),
        .O(\r_xf[7]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBB88888BB88BB8)) 
    \r_xf[7]_i_2 
       (.I0(o_text_out[7]),
        .I1(w_wf_post_pre),
        .I2(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]15_out [7]),
        .I3(o_text_out[63]),
        .I4(\w_rf_mv[0]0 [7]),
        .I5(i_op),
        .O(\r_xf[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_xf[7]_i_4 
       (.I0(i_op),
        .I1(w_rnd_key[6]),
        .O(\r_xf[7]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_xf[7]_i_5 
       (.I0(i_op),
        .I1(w_rnd_key[5]),
        .O(\r_xf[7]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_xf[7]_i_6 
       (.I0(i_op),
        .I1(w_rnd_key[4]),
        .O(\r_xf[7]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBF80407F407FBF80)) 
    \r_xf[7]_i_7 
       (.I0(i_text_in[7]),
        .I1(i_text_val),
        .I2(o_rdy_INST_0_i_1_n_0),
        .I3(o_text_out[7]),
        .I4(w_rnd_key[7]),
        .I5(i_op),
        .O(\r_xf[7]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9699999996666666)) 
    \r_xf[7]_i_8 
       (.I0(w_rnd_key[6]),
        .I1(i_op),
        .I2(i_text_in[6]),
        .I3(i_text_val),
        .I4(o_rdy_INST_0_i_1_n_0),
        .I5(o_text_out[6]),
        .O(\r_xf[7]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9699999996666666)) 
    \r_xf[7]_i_9 
       (.I0(w_rnd_key[5]),
        .I1(i_op),
        .I2(i_text_in[5]),
        .I3(i_text_val),
        .I4(o_rdy_INST_0_i_1_n_0),
        .I5(o_text_out[5]),
        .O(\r_xf[7]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[8]_i_1 
       (.I0(\r_xf[8]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[8]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[8]),
        .O(p_1_in[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \r_xf[8]_i_2 
       (.I0(\w_rf_mv[0]00_in [0]),
        .I1(\w_rf_mv[0]0 [0]),
        .I2(w_wf_post_pre),
        .I3(o_text_out[16]),
        .I4(i_op),
        .I5(o_text_out[0]),
        .O(\r_xf[8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888B8B8B8)) 
    \r_xf[9]_i_1 
       (.I0(\r_xf[9]_i_2_n_0 ),
        .I1(\r_xf[63]_i_9_n_0 ),
        .I2(o_text_out[9]),
        .I3(o_rdy_INST_0_i_1_n_0),
        .I4(i_text_val),
        .I5(i_text_in[9]),
        .O(p_1_in[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \r_xf[9]_i_2 
       (.I0(\w_rf_mv[0]00_in [1]),
        .I1(\w_rf_mv[0]0 [1]),
        .I2(w_wf_post_pre),
        .I3(o_text_out[17]),
        .I4(i_op),
        .I5(o_text_out[1]),
        .O(\r_xf[9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_xf_reg[35]_i_3 
       (.CI(\<const0>__0__0 ),
        .CO(r_xf_reg),
        .CYINIT(\u_CRYPTO_PATH/w_wf_in_mux [32]),
        .DI({\r_xf[35]_i_5_n_0 ,\r_xf[35]_i_6_n_0 ,\r_xf[35]_i_7_n_0 ,i_op}),
        .O({\r_xf_reg[35]_i_3_n_4 ,\r_xf_reg[35]_i_3_n_5 ,\r_xf_reg[35]_i_3_n_6 ,\r_xf_reg[35]_i_3_n_7 }),
        .S({\r_xf[35]_i_8_n_0 ,\r_xf[35]_i_9_n_0 ,\r_xf[35]_i_10_n_0 ,w_rnd_key[16]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_xf_reg[39]_i_3 
       (.CI(r_xf_reg[3]),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\r_xf[39]_i_4_n_0 ,\r_xf[39]_i_5_n_0 ,\r_xf[39]_i_6_n_0 }),
        .O({\r_xf_reg[39]_i_3_n_4 ,\r_xf_reg[39]_i_3_n_5 ,\r_xf_reg[39]_i_3_n_6 ,\r_xf_reg[39]_i_3_n_7 }),
        .S({\r_xf[39]_i_7_n_0 ,\r_xf[39]_i_8_n_0 ,\r_xf[39]_i_9_n_0 ,\r_xf[39]_i_10_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_xf_reg[3]_i_3 
       (.CI(\<const0>__0__0 ),
        .CO({\r_xf_reg[3]_i_3_n_0 ,\r_xf_reg[3]_i_3_n_1 ,\r_xf_reg[3]_i_3_n_2 ,\r_xf_reg[3]_i_3_n_3 }),
        .CYINIT(\u_CRYPTO_PATH/w_wf_in_mux [0]),
        .DI({\r_xf[3]_i_5_n_0 ,\r_xf[3]_i_6_n_0 ,\r_xf[3]_i_7_n_0 ,i_op}),
        .O({\r_xf_reg[3]_i_3_n_4 ,\r_xf_reg[3]_i_3_n_5 ,\r_xf_reg[3]_i_3_n_6 ,\r_xf_reg[3]_i_3_n_7 }),
        .S({\r_xf[3]_i_8_n_0 ,\r_xf[3]_i_9_n_0 ,\r_xf[3]_i_10_n_0 ,w_rnd_key[0]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_xf_reg[7]_i_3 
       (.CI(\r_xf_reg[3]_i_3_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\r_xf[7]_i_4_n_0 ,\r_xf[7]_i_5_n_0 ,\r_xf[7]_i_6_n_0 }),
        .O({\r_xf_reg[7]_i_3_n_4 ,\r_xf_reg[7]_i_3_n_5 ,\r_xf_reg[7]_i_3_n_6 ,\r_xf_reg[7]_i_3_n_7 }),
        .S({\r_xf[7]_i_7_n_0 ,\r_xf[7]_i_8_n_0 ,\r_xf[7]_i_9_n_0 ,\r_xf[7]_i_10_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \u_CONTROL/FSM_sequential_r_pstate_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(FSM_sequential_r_pstate),
        .PRE(\r_xf[63]_i_3_n_0 ),
        .Q(\u_CONTROL/r_pstate [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CONTROL/FSM_sequential_r_pstate_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\FSM_sequential_r_pstate[1]_i_1_n_0 ),
        .Q(\u_CONTROL/r_pstate [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CONTROL/FSM_sequential_r_pstate_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\FSM_sequential_r_pstate[2]_i_1_n_0 ),
        .Q(\u_CONTROL/r_pstate [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CONTROL/FSM_sequential_r_pstate_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\FSM_sequential_r_pstate[3]_i_1_n_0 ),
        .Q(\u_CONTROL/r_pstate [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CONTROL/FSM_sequential_r_pstate_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\FSM_sequential_r_pstate[4]_i_1_n_0 ),
        .Q(\u_CONTROL/r_pstate [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CONTROL/FSM_sequential_r_pstate_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\FSM_sequential_r_pstate[5]_i_1_n_0 ),
        .Q(\u_CONTROL/r_pstate [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[0] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[0]),
        .Q(o_text_out[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[10] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[10]),
        .Q(o_text_out[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[11] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[11]),
        .Q(o_text_out[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[12] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[12]),
        .Q(o_text_out[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[13] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[13]),
        .Q(o_text_out[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[14] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[14]),
        .Q(o_text_out[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[15] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[15]),
        .Q(o_text_out[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[16] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[16]),
        .Q(o_text_out[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[17] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[17]),
        .Q(o_text_out[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[18] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[18]),
        .Q(o_text_out[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[19] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[19]),
        .Q(o_text_out[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[1] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[1]),
        .Q(o_text_out[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[20] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[20]),
        .Q(o_text_out[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[21] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[21]),
        .Q(o_text_out[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[22] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[22]),
        .Q(o_text_out[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[23] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[23]),
        .Q(o_text_out[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[24] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[24]),
        .Q(o_text_out[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[25] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[25]),
        .Q(o_text_out[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[26] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[26]),
        .Q(o_text_out[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[27] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[27]),
        .Q(o_text_out[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[28] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[28]),
        .Q(o_text_out[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[29] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[29]),
        .Q(o_text_out[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[2] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[2]),
        .Q(o_text_out[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[30] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[30]),
        .Q(o_text_out[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[31] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[31]),
        .Q(o_text_out[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[32] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[32]),
        .Q(o_text_out[32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[33] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[33]),
        .Q(o_text_out[33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[34] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[34]),
        .Q(o_text_out[34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[35] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[35]),
        .Q(o_text_out[35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[36] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[36]),
        .Q(o_text_out[36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[37] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[37]),
        .Q(o_text_out[37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[38] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[38]),
        .Q(o_text_out[38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[39] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[39]),
        .Q(o_text_out[39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[3] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[3]),
        .Q(o_text_out[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[40] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[40]),
        .Q(o_text_out[40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[41] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[41]),
        .Q(o_text_out[41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[42] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[42]),
        .Q(o_text_out[42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[43] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[43]),
        .Q(o_text_out[43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[44] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[44]),
        .Q(o_text_out[44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[45] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[45]),
        .Q(o_text_out[45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[46] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[46]),
        .Q(o_text_out[46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[47] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[47]),
        .Q(o_text_out[47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[48] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[48]),
        .Q(o_text_out[48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[49] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[49]),
        .Q(o_text_out[49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[4] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[4]),
        .Q(o_text_out[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[50] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[50]),
        .Q(o_text_out[50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[51] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[51]),
        .Q(o_text_out[51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[52] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[52]),
        .Q(o_text_out[52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[53] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[53]),
        .Q(o_text_out[53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[54] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[54]),
        .Q(o_text_out[54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[55] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[55]),
        .Q(o_text_out[55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[56] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[56]),
        .Q(o_text_out[56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[57] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[57]),
        .Q(o_text_out[57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[58] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[58]),
        .Q(o_text_out[58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[59] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[59]),
        .Q(o_text_out[59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[5] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[5]),
        .Q(o_text_out[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[60] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[60]),
        .Q(o_text_out[60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[61] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[61]),
        .Q(o_text_out[61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[62] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[62]),
        .Q(o_text_out[62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[63] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[63]),
        .Q(o_text_out[63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[6] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[6]),
        .Q(o_text_out[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[7] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[7]),
        .Q(o_text_out[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[8] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[8]),
        .Q(o_text_out[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_CRYPTO_PATH/r_xf_reg[9] 
       (.C(clk),
        .CE(\r_xf[63]_i_1_n_0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_1_in[9]),
        .Q(o_text_out[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_CRYPTO_PATH/u_RF/w_rf_mv[0]0__21_carry 
       (.CI(\<const0>__0__0 ),
        .CO(\u_CRYPTO_PATH/u_RF/w_rf_mv ),
        .CYINIT(\<const0>__0__0 ),
        .DI(o_text_out[11:8]),
        .O(\w_rf_mv[0]00_in [3:0]),
        .S({\w_rf_mv[0]0__21_carry_i_1_n_0 ,\w_rf_mv[0]0__21_carry_i_2_n_0 ,\w_rf_mv[0]0__21_carry_i_3_n_0 ,\w_rf_mv[0]0__21_carry_i_4_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_CRYPTO_PATH/u_RF/w_rf_mv[0]0__21_carry__0 
       (.CI(\u_CRYPTO_PATH/u_RF/w_rf_mv [3]),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,o_text_out[14:12]}),
        .O(\w_rf_mv[0]00_in [7:4]),
        .S({w_rf_mv,\w_rf_mv[0]0__21_carry__0_i_2_n_0 ,\w_rf_mv[0]0__21_carry__0_i_3_n_0 ,\w_rf_mv[0]0__21_carry__0_i_4_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_CRYPTO_PATH/u_RF/w_rf_mv[0]0_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_CRYPTO_PATH/u_RF/w_rf_mv[0]0_carry_n_0 ,\u_CRYPTO_PATH/u_RF/w_rf_mv[0]0_carry_n_1 ,\u_CRYPTO_PATH/u_RF/w_rf_mv[0]0_carry_n_2 ,\u_CRYPTO_PATH/u_RF/w_rf_mv[0]0_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI(o_text_out[11:8]),
        .O(\w_rf_mv[0]0 [3:0]),
        .S({\w_rf_mv[0]0_carry_i_1_n_0 ,\w_rf_mv[0]0_carry_i_2_n_0 ,\w_rf_mv[0]0_carry_i_3_n_0 ,\w_rf_mv[0]0_carry_i_4_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_CRYPTO_PATH/u_RF/w_rf_mv[0]0_carry__0 
       (.CI(\u_CRYPTO_PATH/u_RF/w_rf_mv[0]0_carry_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,o_text_out[14:12]}),
        .O(\w_rf_mv[0]0 [7:4]),
        .S({\w_rf_mv[0]0_carry__0_i_1_n_0 ,\w_rf_mv[0]0_carry__0_i_2_n_0 ,\w_rf_mv[0]0_carry__0_i_3_n_0 ,\w_rf_mv[0]0_carry__0_i_4_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__21_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__21_carry_n_0 ,\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__21_carry_n_1 ,\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__21_carry_n_2 ,\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__21_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(w_rnd_key[11:8]),
        .O(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]12_out [3:0]),
        .S({\w_rf_mv[1]1__21_carry_i_1_n_0 ,\w_rf_mv[1]1__21_carry_i_2_n_0 ,\w_rf_mv[1]1__21_carry_i_3_n_0 ,\w_rf_mv[1]1__21_carry_i_4_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__21_carry__0 
       (.CI(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__21_carry_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,w_rnd_key[14:12]}),
        .O(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]12_out [7:4]),
        .S({\w_rf_mv[1]1__21_carry__0_i_1_n_0 ,\w_rf_mv[1]1__21_carry__0_i_2_n_0 ,\w_rf_mv[1]1__21_carry__0_i_3_n_0 ,\w_rf_mv[1]1__21_carry__0_i_4_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_CRYPTO_PATH/u_RF/w_rf_mv[1]1_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1_carry_n_0 ,\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1_carry_n_1 ,\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1_carry_n_2 ,\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(w_rnd_key[19:16]),
        .O(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__43 [3:0]),
        .S({\w_rf_mv[1]1_carry_i_1_n_0 ,\w_rf_mv[1]1_carry_i_2_n_0 ,\w_rf_mv[1]1_carry_i_3_n_0 ,\w_rf_mv[1]1_carry_i_4_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_CRYPTO_PATH/u_RF/w_rf_mv[1]1_carry__0 
       (.CI(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1_carry_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,w_rnd_key[22:20]}),
        .O(\u_CRYPTO_PATH/u_RF/w_rf_mv[1]1__43 [7:4]),
        .S({\w_rf_mv[1]1_carry__0_i_1_n_0 ,\w_rf_mv[1]1_carry__0_i_2_n_0 ,\w_rf_mv[1]1_carry__0_i_3_n_0 ,\w_rf_mv[1]1_carry__0_i_4_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_CRYPTO_PATH/u_RF/w_rf_mv[2]0__21_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_CRYPTO_PATH/u_RF/w_rf_mv[2]0__21_carry_n_0 ,\u_CRYPTO_PATH/u_RF/w_rf_mv[2]0__21_carry_n_1 ,\u_CRYPTO_PATH/u_RF/w_rf_mv[2]0__21_carry_n_2 ,\u_CRYPTO_PATH/u_RF/w_rf_mv[2]0__21_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(o_text_out[43:40]),
        .O(\w_rf_mv[2]01_in [3:0]),
        .S({\w_rf_mv[2]0__21_carry_i_1_n_0 ,\w_rf_mv[2]0__21_carry_i_2_n_0 ,\w_rf_mv[2]0__21_carry_i_3_n_0 ,\w_rf_mv[2]0__21_carry_i_4_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_CRYPTO_PATH/u_RF/w_rf_mv[2]0__21_carry__0 
       (.CI(\u_CRYPTO_PATH/u_RF/w_rf_mv[2]0__21_carry_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,o_text_out[46:44]}),
        .O(\w_rf_mv[2]01_in [7:4]),
        .S({\w_rf_mv[2]0__21_carry__0_i_1_n_0 ,\w_rf_mv[2]0__21_carry__0_i_2_n_0 ,\w_rf_mv[2]0__21_carry__0_i_3_n_0 ,\w_rf_mv[2]0__21_carry__0_i_4_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_CRYPTO_PATH/u_RF/w_rf_mv[2]0_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_CRYPTO_PATH/u_RF/w_rf_mv[2]0_carry_n_0 ,\u_CRYPTO_PATH/u_RF/w_rf_mv[2]0_carry_n_1 ,\u_CRYPTO_PATH/u_RF/w_rf_mv[2]0_carry_n_2 ,\u_CRYPTO_PATH/u_RF/w_rf_mv[2]0_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI(o_text_out[43:40]),
        .O(\w_rf_mv[2]0 [3:0]),
        .S({\w_rf_mv[2]0_carry_i_1_n_0 ,\w_rf_mv[2]0_carry_i_2_n_0 ,\w_rf_mv[2]0_carry_i_3_n_0 ,\w_rf_mv[2]0_carry_i_4_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_CRYPTO_PATH/u_RF/w_rf_mv[2]0_carry__0 
       (.CI(\u_CRYPTO_PATH/u_RF/w_rf_mv[2]0_carry_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,o_text_out[46:44]}),
        .O(\w_rf_mv[2]0 [7:4]),
        .S({\w_rf_mv[2]0_carry__0_i_1_n_0 ,\w_rf_mv[2]0_carry__0_i_2_n_0 ,\w_rf_mv[2]0_carry__0_i_3_n_0 ,\w_rf_mv[2]0_carry__0_i_4_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__21_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__21_carry_n_0 ,\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__21_carry_n_1 ,\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__21_carry_n_2 ,\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__21_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(w_rnd_key[3:0]),
        .O(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__43 [3:0]),
        .S({\w_rf_mv[3]1__21_carry_i_1__0_n_0 ,\w_rf_mv[3]1__21_carry_i_2_n_0 ,\w_rf_mv[3]1__21_carry_i_3_n_0 ,\w_rf_mv[3]1__21_carry_i_4_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__21_carry__0 
       (.CI(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__21_carry_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,w_rnd_key[6:4]}),
        .O(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1__43 [7:4]),
        .S({\w_rf_mv[3]1__21_carry_i_1_n_0 ,\w_rf_mv[3]1__21_carry_i_2__0_n_0 ,\w_rf_mv[3]1__21_carry_i_3__0_n_0 ,\w_rf_mv[3]1__21_carry_i_4__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_CRYPTO_PATH/u_RF/w_rf_mv[3]1_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1_carry_n_0 ,\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1_carry_n_1 ,\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1_carry_n_2 ,\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(w_rnd_key[27:24]),
        .O(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]15_out [3:0]),
        .S({\w_rf_mv[3]1_carry_i_1_n_0 ,\w_rf_mv[3]1_carry_i_2_n_0 ,\w_rf_mv[3]1_carry_i_3_n_0 ,\w_rf_mv[3]1_carry_i_4_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_CRYPTO_PATH/u_RF/w_rf_mv[3]1_carry__0 
       (.CI(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]1_carry_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,w_rnd_key[30:28]}),
        .O(\u_CRYPTO_PATH/u_RF/w_rf_mv[3]15_out [7:4]),
        .S({\w_rf_mv[3]1_carry__0_i_1_n_0 ,\w_rf_mv[3]1_carry__0_i_2_n_0 ,\w_rf_mv[3]1_carry__0_i_3_n_0 ,\w_rf_mv[3]1_carry__0_i_4_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_0x_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_0_in[0]),
        .Q(w_rnd_key[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_0x_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_0_in[1]),
        .Q(w_rnd_key[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_0x_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_0_in[2]),
        .Q(w_rnd_key[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_0x_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_0_in[3]),
        .Q(w_rnd_key[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_0x_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_0_in[4]),
        .Q(w_rnd_key[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_0x_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_0_in[5]),
        .Q(w_rnd_key[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_0x_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_0_in[6]),
        .Q(w_rnd_key[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_0x_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(p_0_in[7]),
        .Q(w_rnd_key[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_1x_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(r_rnd_key_1x),
        .Q(w_rnd_key[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_1x_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\r_rnd_key_1x[1]_i_1_n_0 ),
        .Q(w_rnd_key[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_1x_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\r_rnd_key_1x[2]_i_1_n_0 ),
        .Q(w_rnd_key[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_1x_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\r_rnd_key_1x[3]_i_1_n_0 ),
        .Q(w_rnd_key[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_1x_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\r_rnd_key_1x[4]_i_1_n_0 ),
        .Q(w_rnd_key[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_1x_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\r_rnd_key_1x[5]_i_1_n_0 ),
        .Q(w_rnd_key[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_1x_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\r_rnd_key_1x[6]_i_1_n_0 ),
        .Q(w_rnd_key[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_1x_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\r_rnd_key_1x[7]_i_1_n_0 ),
        .Q(w_rnd_key[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_2x_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(r_rnd_key_2x),
        .Q(w_rnd_key[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_2x_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\r_rnd_key_2x[1]_i_1_n_0 ),
        .Q(w_rnd_key[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_2x_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\r_rnd_key_2x[2]_i_1_n_0 ),
        .Q(w_rnd_key[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_2x_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\r_rnd_key_2x[3]_i_1_n_0 ),
        .Q(w_rnd_key[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_2x_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\r_rnd_key_2x[4]_i_1_n_0 ),
        .Q(w_rnd_key[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_2x_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\r_rnd_key_2x[5]_i_1_n_0 ),
        .Q(w_rnd_key[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_2x_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\r_rnd_key_2x[6]_i_1_n_0 ),
        .Q(w_rnd_key[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_2x_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\r_rnd_key_2x[7]_i_1_n_0 ),
        .Q(w_rnd_key[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_3x_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(r_rnd_key_3x),
        .Q(w_rnd_key[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_3x_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\r_rnd_key_3x[1]_i_1_n_0 ),
        .Q(w_rnd_key[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_3x_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\r_rnd_key_3x[2]_i_1_n_0 ),
        .Q(w_rnd_key[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_3x_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\r_rnd_key_3x[3]_i_1_n_0 ),
        .Q(w_rnd_key[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_3x_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\r_rnd_key_3x[4]_i_1_n_0 ),
        .Q(w_rnd_key[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_3x_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\r_rnd_key_3x[5]_i_1_n_0 ),
        .Q(w_rnd_key[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_3x_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\r_rnd_key_3x[6]_i_1_n_0 ),
        .Q(w_rnd_key[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \u_KEY_SCHED/r_rnd_key_3x_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\r_xf[63]_i_3_n_0 ),
        .D(\r_rnd_key_3x[7]_i_1_n_0 ),
        .Q(w_rnd_key[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_10 
       (.I0(g0_b2_n_0),
        .I1(\r_rnd_key_0x[3]_i_28_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[3]_i_29_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[3]_i_30_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_0x ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_11 
       (.I0(g0_b1_n_0),
        .I1(\r_rnd_key_0x[3]_i_31_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[3]_i_32_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[3]_i_33_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_12 
       (.I0(g0_b0_n_0),
        .I1(\r_rnd_key_0x[3]_i_34_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[3]_i_35_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[3]_i_36_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_5 
       (.I0(g0_b6_n_0),
        .I1(\r_rnd_key_0x[3]_i_13_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[3]_i_14_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[3]_i_15_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_6 
       (.I0(g0_b5_n_0),
        .I1(\r_rnd_key_0x[3]_i_16_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[3]_i_17_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[3]_i_18_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_7 
       (.I0(g0_b4_n_0),
        .I1(\r_rnd_key_0x[3]_i_19_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[3]_i_20_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[3]_i_21_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_8 
       (.I0(g0_b0__0_n_0),
        .I1(\r_rnd_key_0x[3]_i_22_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[3]_i_23_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[3]_i_24_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_9 
       (.I0(g0_b0__0_n_0),
        .I1(\r_rnd_key_0x[3]_i_25_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[3]_i_26_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[3]_i_27_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_0x[3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_0x[7]_i_11 
       (.I0(g0_b6_n_0),
        .I1(\r_rnd_key_0x[7]_i_31_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[7]_i_32_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[7]_i_33_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_0x[7]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_0x[7]_i_12 
       (.I0(g0_b5_n_0),
        .I1(\r_rnd_key_0x[7]_i_34_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[7]_i_35_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[7]_i_36_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_0x[7]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_0x[7]_i_13 
       (.I0(g0_b4_n_0),
        .I1(\r_rnd_key_0x[7]_i_37_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[7]_i_38_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[7]_i_39_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_0x[7]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_0x[7]_i_7 
       (.I0(g0_b6__0_n_0),
        .I1(\r_rnd_key_0x[7]_i_18_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[7]_i_19_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[7]_i_20_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_0x[7]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_0x[7]_i_8 
       (.I0(g0_b5__0_n_0),
        .I1(\r_rnd_key_0x[7]_i_21_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[7]_i_22_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[7]_i_23_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_0x[7]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_0x[7]_i_9 
       (.I0(g0_b4__0_n_0),
        .I1(\r_rnd_key_0x[7]_i_24_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[7]_i_25_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[7]_i_26_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_0x[7]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_10 
       (.I0(g0_b0__0_n_0),
        .I1(\r_rnd_key_1x[3]_i_23_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[3]_i_18_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_1x[3]_i_24_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_1x ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_11 
       (.I0(g0_b2_n_0),
        .I1(\r_rnd_key_1x[3]_i_25_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[3]_i_21_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_1x[3]_i_26_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_12 
       (.I0(g0_b1_n_0),
        .I1(\r_rnd_key_1x[3]_i_27_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[3]_i_24_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_1x[3]_i_28_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_5 
       (.I0(g0_b5_n_0),
        .I1(\r_rnd_key_1x[3]_i_13_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_1x[3]_i_14_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[3]_i_26_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_6 
       (.I0(g0_b4_n_0),
        .I1(\r_rnd_key_1x[3]_i_15_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_1x[3]_i_16_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[3]_i_29_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_7 
       (.I0(g0_b0__0_n_0),
        .I1(\r_rnd_key_1x[3]_i_17_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_1x[3]_i_18_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[3]_i_32_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_8 
       (.I0(g0_b2_n_0),
        .I1(\r_rnd_key_1x[3]_i_19_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_1x[3]_i_20_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[3]_i_35_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_9 
       (.I0(g0_b4_n_0),
        .I1(\r_rnd_key_1x[3]_i_21_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[3]_i_15_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_1x[3]_i_22_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_1x[3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_1x[7]_i_10 
       (.I0(g0_b4__0_n_0),
        .I1(\r_rnd_key_1x[7]_i_19_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[7]_i_20_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_1x[7]_i_20_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_1x[7]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_1x[7]_i_11 
       (.I0(g0_b6_n_0),
        .I1(\r_rnd_key_1x[7]_i_21_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[7]_i_23_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_1x[7]_i_22_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_1x[7]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_1x[7]_i_12 
       (.I0(g0_b5_n_0),
        .I1(\r_rnd_key_1x[7]_i_23_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_0x[7]_i_26_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_1x[7]_i_24_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_1x[7]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_1x[7]_i_6 
       (.I0(g0_b5__0_n_0),
        .I1(\r_rnd_key_1x[7]_i_13_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_1x[7]_i_14_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[7]_i_32_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_1x[7]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_1x[7]_i_7 
       (.I0(g0_b4__0_n_0),
        .I1(\r_rnd_key_1x[7]_i_15_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_1x[7]_i_16_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[7]_i_35_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_1x[7]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h565656A6A6A656A6)) 
    \u_KEY_SCHED/u_SKG/r_rnd_key_1x[7]_i_8 
       (.I0(g0_b6_n_0),
        .I1(\r_rnd_key_1x[7]_i_17_n_0 ),
        .I2(\u_KEY_SCHED/u_SKG/w_base [4]),
        .I3(\r_rnd_key_1x[7]_i_18_n_0 ),
        .I4(\u_KEY_SCHED/u_SKG/w_base [3]),
        .I5(\r_rnd_key_0x[7]_i_38_n_0 ),
        .O(\u_KEY_SCHED/u_SKG/r_rnd_key_1x[7]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \w_rf_mv[0]0__21_carry__0_i_1 
       (.I0(o_text_out[3]),
        .I1(o_text_out[4]),
        .I2(o_text_out[1]),
        .I3(w_rnd_key[7]),
        .I4(o_text_out[15]),
        .O(w_rf_mv));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \w_rf_mv[0]0__21_carry__0_i_2 
       (.I0(o_text_out[14]),
        .I1(o_text_out[0]),
        .I2(o_text_out[3]),
        .I3(o_text_out[2]),
        .I4(w_rnd_key[6]),
        .O(\w_rf_mv[0]0__21_carry__0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \w_rf_mv[0]0__21_carry__0_i_3 
       (.I0(o_text_out[13]),
        .I1(o_text_out[1]),
        .I2(o_text_out[7]),
        .I3(o_text_out[2]),
        .I4(w_rnd_key[5]),
        .O(\w_rf_mv[0]0__21_carry__0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \w_rf_mv[0]0__21_carry__0_i_4 
       (.I0(o_text_out[12]),
        .I1(o_text_out[0]),
        .I2(o_text_out[6]),
        .I3(o_text_out[1]),
        .I4(w_rnd_key[4]),
        .O(\w_rf_mv[0]0__21_carry__0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \w_rf_mv[0]0__21_carry_i_1 
       (.I0(o_text_out[11]),
        .I1(o_text_out[0]),
        .I2(o_text_out[7]),
        .I3(o_text_out[5]),
        .I4(w_rnd_key[3]),
        .O(\w_rf_mv[0]0__21_carry_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \w_rf_mv[0]0__21_carry_i_2 
       (.I0(o_text_out[10]),
        .I1(o_text_out[4]),
        .I2(o_text_out[7]),
        .I3(o_text_out[6]),
        .I4(w_rnd_key[2]),
        .O(\w_rf_mv[0]0__21_carry_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \w_rf_mv[0]0__21_carry_i_3 
       (.I0(o_text_out[9]),
        .I1(o_text_out[3]),
        .I2(o_text_out[6]),
        .I3(o_text_out[5]),
        .I4(w_rnd_key[1]),
        .O(\w_rf_mv[0]0__21_carry_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \w_rf_mv[0]0__21_carry_i_4 
       (.I0(o_text_out[8]),
        .I1(o_text_out[2]),
        .I2(o_text_out[5]),
        .I3(o_text_out[4]),
        .I4(w_rnd_key[0]),
        .O(\w_rf_mv[0]0__21_carry_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969669)) 
    \w_rf_mv[0]0_carry__0_i_1 
       (.I0(o_text_out[3]),
        .I1(o_text_out[4]),
        .I2(o_text_out[1]),
        .I3(w_rnd_key[31]),
        .I4(o_text_out[15]),
        .O(\w_rf_mv[0]0_carry__0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969669)) 
    \w_rf_mv[0]0_carry__0_i_2 
       (.I0(o_text_out[14]),
        .I1(o_text_out[0]),
        .I2(o_text_out[3]),
        .I3(o_text_out[2]),
        .I4(w_rnd_key[30]),
        .O(\w_rf_mv[0]0_carry__0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969669)) 
    \w_rf_mv[0]0_carry__0_i_3 
       (.I0(o_text_out[13]),
        .I1(o_text_out[1]),
        .I2(o_text_out[7]),
        .I3(o_text_out[2]),
        .I4(w_rnd_key[29]),
        .O(\w_rf_mv[0]0_carry__0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969669)) 
    \w_rf_mv[0]0_carry__0_i_4 
       (.I0(o_text_out[12]),
        .I1(o_text_out[0]),
        .I2(o_text_out[6]),
        .I3(o_text_out[1]),
        .I4(w_rnd_key[28]),
        .O(\w_rf_mv[0]0_carry__0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969669)) 
    \w_rf_mv[0]0_carry_i_1 
       (.I0(o_text_out[11]),
        .I1(o_text_out[0]),
        .I2(o_text_out[7]),
        .I3(o_text_out[5]),
        .I4(w_rnd_key[27]),
        .O(\w_rf_mv[0]0_carry_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969669)) 
    \w_rf_mv[0]0_carry_i_2 
       (.I0(o_text_out[10]),
        .I1(o_text_out[4]),
        .I2(o_text_out[7]),
        .I3(o_text_out[6]),
        .I4(w_rnd_key[26]),
        .O(\w_rf_mv[0]0_carry_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969669)) 
    \w_rf_mv[0]0_carry_i_3 
       (.I0(o_text_out[9]),
        .I1(o_text_out[3]),
        .I2(o_text_out[6]),
        .I3(o_text_out[5]),
        .I4(w_rnd_key[25]),
        .O(\w_rf_mv[0]0_carry_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969669)) 
    \w_rf_mv[0]0_carry_i_4 
       (.I0(o_text_out[8]),
        .I1(o_text_out[2]),
        .I2(o_text_out[5]),
        .I3(o_text_out[4]),
        .I4(w_rnd_key[24]),
        .O(\w_rf_mv[0]0_carry_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[1]1__21_carry__0_i_1 
       (.I0(w_rnd_key[15]),
        .I1(o_text_out[16]),
        .I2(o_text_out[21]),
        .I3(o_text_out[22]),
        .O(\w_rf_mv[1]1__21_carry__0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[1]1__21_carry__0_i_2 
       (.I0(o_text_out[23]),
        .I1(o_text_out[20]),
        .I2(o_text_out[21]),
        .I3(w_rnd_key[14]),
        .O(\w_rf_mv[1]1__21_carry__0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[1]1__21_carry__0_i_3 
       (.I0(o_text_out[22]),
        .I1(o_text_out[19]),
        .I2(o_text_out[20]),
        .I3(w_rnd_key[13]),
        .O(\w_rf_mv[1]1__21_carry__0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[1]1__21_carry__0_i_4 
       (.I0(o_text_out[18]),
        .I1(o_text_out[21]),
        .I2(o_text_out[19]),
        .I3(w_rnd_key[12]),
        .O(\w_rf_mv[1]1__21_carry__0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[1]1__21_carry_i_1 
       (.I0(o_text_out[17]),
        .I1(o_text_out[20]),
        .I2(o_text_out[18]),
        .I3(w_rnd_key[11]),
        .O(\w_rf_mv[1]1__21_carry_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[1]1__21_carry_i_2 
       (.I0(o_text_out[16]),
        .I1(o_text_out[19]),
        .I2(o_text_out[17]),
        .I3(w_rnd_key[10]),
        .O(\w_rf_mv[1]1__21_carry_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[1]1__21_carry_i_3 
       (.I0(o_text_out[23]),
        .I1(o_text_out[18]),
        .I2(o_text_out[16]),
        .I3(w_rnd_key[9]),
        .O(\w_rf_mv[1]1__21_carry_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[1]1__21_carry_i_4 
       (.I0(o_text_out[22]),
        .I1(o_text_out[17]),
        .I2(o_text_out[23]),
        .I3(w_rnd_key[8]),
        .O(\w_rf_mv[1]1__21_carry_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[1]1_carry__0_i_1 
       (.I0(w_rnd_key[23]),
        .I1(o_text_out[16]),
        .I2(o_text_out[21]),
        .I3(o_text_out[22]),
        .O(\w_rf_mv[1]1_carry__0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[1]1_carry__0_i_2 
       (.I0(o_text_out[23]),
        .I1(o_text_out[20]),
        .I2(o_text_out[21]),
        .I3(w_rnd_key[22]),
        .O(\w_rf_mv[1]1_carry__0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[1]1_carry__0_i_3 
       (.I0(o_text_out[22]),
        .I1(o_text_out[19]),
        .I2(o_text_out[20]),
        .I3(w_rnd_key[21]),
        .O(\w_rf_mv[1]1_carry__0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[1]1_carry__0_i_4 
       (.I0(o_text_out[18]),
        .I1(o_text_out[21]),
        .I2(o_text_out[19]),
        .I3(w_rnd_key[20]),
        .O(\w_rf_mv[1]1_carry__0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[1]1_carry_i_1 
       (.I0(o_text_out[17]),
        .I1(o_text_out[20]),
        .I2(o_text_out[18]),
        .I3(w_rnd_key[19]),
        .O(\w_rf_mv[1]1_carry_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[1]1_carry_i_2 
       (.I0(o_text_out[16]),
        .I1(o_text_out[19]),
        .I2(o_text_out[17]),
        .I3(w_rnd_key[18]),
        .O(\w_rf_mv[1]1_carry_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[1]1_carry_i_3 
       (.I0(o_text_out[23]),
        .I1(o_text_out[18]),
        .I2(o_text_out[16]),
        .I3(w_rnd_key[17]),
        .O(\w_rf_mv[1]1_carry_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[1]1_carry_i_4 
       (.I0(o_text_out[22]),
        .I1(o_text_out[17]),
        .I2(o_text_out[23]),
        .I3(w_rnd_key[16]),
        .O(\w_rf_mv[1]1_carry_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \w_rf_mv[2]0__21_carry__0_i_1 
       (.I0(o_text_out[35]),
        .I1(o_text_out[33]),
        .I2(o_text_out[36]),
        .I3(w_rnd_key[23]),
        .I4(o_text_out[47]),
        .O(\w_rf_mv[2]0__21_carry__0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \w_rf_mv[2]0__21_carry__0_i_2 
       (.I0(o_text_out[46]),
        .I1(o_text_out[34]),
        .I2(o_text_out[32]),
        .I3(o_text_out[35]),
        .I4(w_rnd_key[22]),
        .O(\w_rf_mv[2]0__21_carry__0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \w_rf_mv[2]0__21_carry__0_i_3 
       (.I0(o_text_out[45]),
        .I1(o_text_out[34]),
        .I2(o_text_out[33]),
        .I3(o_text_out[39]),
        .I4(w_rnd_key[21]),
        .O(\w_rf_mv[2]0__21_carry__0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \w_rf_mv[2]0__21_carry__0_i_4 
       (.I0(o_text_out[44]),
        .I1(o_text_out[38]),
        .I2(o_text_out[33]),
        .I3(o_text_out[32]),
        .I4(w_rnd_key[20]),
        .O(\w_rf_mv[2]0__21_carry__0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \w_rf_mv[2]0__21_carry_i_1 
       (.I0(o_text_out[43]),
        .I1(o_text_out[37]),
        .I2(o_text_out[32]),
        .I3(o_text_out[39]),
        .I4(w_rnd_key[19]),
        .O(\w_rf_mv[2]0__21_carry_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \w_rf_mv[2]0__21_carry_i_2 
       (.I0(o_text_out[42]),
        .I1(o_text_out[36]),
        .I2(o_text_out[39]),
        .I3(o_text_out[38]),
        .I4(w_rnd_key[18]),
        .O(\w_rf_mv[2]0__21_carry_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \w_rf_mv[2]0__21_carry_i_3 
       (.I0(o_text_out[41]),
        .I1(o_text_out[37]),
        .I2(o_text_out[38]),
        .I3(o_text_out[35]),
        .I4(w_rnd_key[17]),
        .O(\w_rf_mv[2]0__21_carry_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \w_rf_mv[2]0__21_carry_i_4 
       (.I0(o_text_out[40]),
        .I1(o_text_out[36]),
        .I2(o_text_out[37]),
        .I3(o_text_out[34]),
        .I4(w_rnd_key[16]),
        .O(\w_rf_mv[2]0__21_carry_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969669)) 
    \w_rf_mv[2]0_carry__0_i_1 
       (.I0(o_text_out[35]),
        .I1(o_text_out[33]),
        .I2(o_text_out[36]),
        .I3(w_rnd_key[15]),
        .I4(o_text_out[47]),
        .O(\w_rf_mv[2]0_carry__0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969669)) 
    \w_rf_mv[2]0_carry__0_i_2 
       (.I0(o_text_out[46]),
        .I1(o_text_out[34]),
        .I2(o_text_out[32]),
        .I3(o_text_out[35]),
        .I4(w_rnd_key[14]),
        .O(\w_rf_mv[2]0_carry__0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969669)) 
    \w_rf_mv[2]0_carry__0_i_3 
       (.I0(o_text_out[45]),
        .I1(o_text_out[34]),
        .I2(o_text_out[33]),
        .I3(o_text_out[39]),
        .I4(w_rnd_key[13]),
        .O(\w_rf_mv[2]0_carry__0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969669)) 
    \w_rf_mv[2]0_carry__0_i_4 
       (.I0(o_text_out[44]),
        .I1(o_text_out[38]),
        .I2(o_text_out[33]),
        .I3(o_text_out[32]),
        .I4(w_rnd_key[12]),
        .O(\w_rf_mv[2]0_carry__0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969669)) 
    \w_rf_mv[2]0_carry_i_1 
       (.I0(o_text_out[43]),
        .I1(o_text_out[37]),
        .I2(o_text_out[32]),
        .I3(o_text_out[39]),
        .I4(w_rnd_key[11]),
        .O(\w_rf_mv[2]0_carry_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969669)) 
    \w_rf_mv[2]0_carry_i_2 
       (.I0(o_text_out[42]),
        .I1(o_text_out[36]),
        .I2(o_text_out[39]),
        .I3(o_text_out[38]),
        .I4(w_rnd_key[10]),
        .O(\w_rf_mv[2]0_carry_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969669)) 
    \w_rf_mv[2]0_carry_i_3 
       (.I0(o_text_out[41]),
        .I1(o_text_out[37]),
        .I2(o_text_out[38]),
        .I3(o_text_out[35]),
        .I4(w_rnd_key[9]),
        .O(\w_rf_mv[2]0_carry_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969669)) 
    \w_rf_mv[2]0_carry_i_4 
       (.I0(o_text_out[40]),
        .I1(o_text_out[36]),
        .I2(o_text_out[37]),
        .I3(o_text_out[34]),
        .I4(w_rnd_key[8]),
        .O(\w_rf_mv[2]0_carry_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[3]1__21_carry_i_1 
       (.I0(w_rnd_key[7]),
        .I1(o_text_out[48]),
        .I2(o_text_out[53]),
        .I3(o_text_out[54]),
        .O(\w_rf_mv[3]1__21_carry_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[3]1__21_carry_i_1__0 
       (.I0(o_text_out[49]),
        .I1(o_text_out[52]),
        .I2(o_text_out[50]),
        .I3(w_rnd_key[3]),
        .O(\w_rf_mv[3]1__21_carry_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[3]1__21_carry_i_2 
       (.I0(o_text_out[48]),
        .I1(o_text_out[51]),
        .I2(o_text_out[49]),
        .I3(w_rnd_key[2]),
        .O(\w_rf_mv[3]1__21_carry_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[3]1__21_carry_i_2__0 
       (.I0(o_text_out[55]),
        .I1(o_text_out[52]),
        .I2(o_text_out[53]),
        .I3(w_rnd_key[6]),
        .O(\w_rf_mv[3]1__21_carry_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[3]1__21_carry_i_3 
       (.I0(o_text_out[55]),
        .I1(o_text_out[50]),
        .I2(o_text_out[48]),
        .I3(w_rnd_key[1]),
        .O(\w_rf_mv[3]1__21_carry_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[3]1__21_carry_i_3__0 
       (.I0(o_text_out[54]),
        .I1(o_text_out[51]),
        .I2(o_text_out[52]),
        .I3(w_rnd_key[5]),
        .O(\w_rf_mv[3]1__21_carry_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[3]1__21_carry_i_4 
       (.I0(o_text_out[54]),
        .I1(o_text_out[49]),
        .I2(o_text_out[55]),
        .I3(w_rnd_key[0]),
        .O(\w_rf_mv[3]1__21_carry_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[3]1__21_carry_i_4__0 
       (.I0(o_text_out[50]),
        .I1(o_text_out[53]),
        .I2(o_text_out[51]),
        .I3(w_rnd_key[4]),
        .O(\w_rf_mv[3]1__21_carry_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[3]1_carry__0_i_1 
       (.I0(w_rnd_key[31]),
        .I1(o_text_out[48]),
        .I2(o_text_out[53]),
        .I3(o_text_out[54]),
        .O(\w_rf_mv[3]1_carry__0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[3]1_carry__0_i_2 
       (.I0(o_text_out[55]),
        .I1(o_text_out[52]),
        .I2(o_text_out[53]),
        .I3(w_rnd_key[30]),
        .O(\w_rf_mv[3]1_carry__0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[3]1_carry__0_i_3 
       (.I0(o_text_out[54]),
        .I1(o_text_out[51]),
        .I2(o_text_out[52]),
        .I3(w_rnd_key[29]),
        .O(\w_rf_mv[3]1_carry__0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[3]1_carry__0_i_4 
       (.I0(o_text_out[50]),
        .I1(o_text_out[53]),
        .I2(o_text_out[51]),
        .I3(w_rnd_key[28]),
        .O(\w_rf_mv[3]1_carry__0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[3]1_carry_i_1 
       (.I0(o_text_out[49]),
        .I1(o_text_out[52]),
        .I2(o_text_out[50]),
        .I3(w_rnd_key[27]),
        .O(\w_rf_mv[3]1_carry_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[3]1_carry_i_2 
       (.I0(o_text_out[48]),
        .I1(o_text_out[51]),
        .I2(o_text_out[49]),
        .I3(w_rnd_key[26]),
        .O(\w_rf_mv[3]1_carry_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[3]1_carry_i_3 
       (.I0(o_text_out[55]),
        .I1(o_text_out[50]),
        .I2(o_text_out[48]),
        .I3(w_rnd_key[25]),
        .O(\w_rf_mv[3]1_carry_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \w_rf_mv[3]1_carry_i_4 
       (.I0(o_text_out[54]),
        .I1(o_text_out[49]),
        .I2(o_text_out[55]),
        .I3(w_rnd_key[24]),
        .O(\w_rf_mv[3]1_carry_i_4_n_0 ));
endmodule
